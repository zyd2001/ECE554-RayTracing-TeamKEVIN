// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.2.0 Build 57 06/24/2019 Patches 0.01dc SJ Pro Edition"

// DATE "04/20/2021 23:13:10"

// 
// Device: Altera 1SX280HN2F43E2VG Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Fix_Div (
	result,
	clk,
	rst,
	en,
	denominator,
	numerator)/* synthesis synthesis_greybox=0 */;
output 	[31:0] result;
input 	clk;
input 	rst;
input 	[0:0] en;
input 	[31:0] denominator;
input 	[31:0] numerator;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a_aq;
wire fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a_aq;
wire fxp_functions_0_aadd_17_a1_sumout;
wire fxp_functions_0_aadd_17_a2;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a_aq;
wire fxp_functions_0_aadd_17_a6_sumout;
wire fxp_functions_0_aadd_17_a7;
wire fxp_functions_0_aadd_17_a11_sumout;
wire fxp_functions_0_aadd_17_a12;
wire fxp_functions_0_aadd_17_a16_sumout;
wire fxp_functions_0_aadd_17_a17;
wire fxp_functions_0_aadd_17_a21_sumout;
wire fxp_functions_0_aadd_17_a22;
wire fxp_functions_0_aadd_17_a26_sumout;
wire fxp_functions_0_aadd_17_a27;
wire fxp_functions_0_aadd_17_a31_sumout;
wire fxp_functions_0_aadd_17_a32;
wire fxp_functions_0_aadd_17_a36_sumout;
wire fxp_functions_0_aadd_17_a37;
wire fxp_functions_0_aadd_17_a41_sumout;
wire fxp_functions_0_aadd_17_a42;
wire fxp_functions_0_aadd_17_a46_sumout;
wire fxp_functions_0_aadd_17_a47;
wire fxp_functions_0_aadd_17_a51_sumout;
wire fxp_functions_0_aadd_17_a52;
wire fxp_functions_0_aadd_17_a56_sumout;
wire fxp_functions_0_aadd_17_a57;
wire fxp_functions_0_aadd_17_a61_sumout;
wire fxp_functions_0_aadd_17_a62;
wire fxp_functions_0_aadd_17_a66_sumout;
wire fxp_functions_0_aadd_17_a67;
wire fxp_functions_0_aadd_17_a71_sumout;
wire fxp_functions_0_aadd_17_a72;
wire fxp_functions_0_aadd_17_a76_sumout;
wire fxp_functions_0_aadd_17_a77;
wire fxp_functions_0_aadd_17_a81_sumout;
wire fxp_functions_0_aadd_17_a82;
wire fxp_functions_0_aadd_17_a86_sumout;
wire fxp_functions_0_aadd_17_a87;
wire fxp_functions_0_aadd_17_a91_sumout;
wire fxp_functions_0_aadd_17_a92;
wire fxp_functions_0_aadd_17_a96_sumout;
wire fxp_functions_0_aadd_17_a97;
wire fxp_functions_0_aadd_17_a101_sumout;
wire fxp_functions_0_aadd_17_a102;
wire fxp_functions_0_aadd_17_a106_sumout;
wire fxp_functions_0_aadd_17_a107;
wire fxp_functions_0_aadd_17_a111_sumout;
wire fxp_functions_0_aadd_17_a112;
wire fxp_functions_0_aadd_17_a116_sumout;
wire fxp_functions_0_aadd_17_a117;
wire fxp_functions_0_aadd_17_a121_sumout;
wire fxp_functions_0_aadd_17_a122;
wire fxp_functions_0_aadd_17_a126_sumout;
wire fxp_functions_0_aadd_17_a127;
wire fxp_functions_0_aadd_17_a131_sumout;
wire fxp_functions_0_aadd_17_a132;
wire fxp_functions_0_aadd_17_a136_sumout;
wire fxp_functions_0_aadd_17_a137;
wire fxp_functions_0_aadd_17_a141_sumout;
wire fxp_functions_0_aadd_17_a142;
wire fxp_functions_0_aadd_17_a146_sumout;
wire fxp_functions_0_aadd_17_a147;
wire fxp_functions_0_aadd_17_a151_sumout;
wire fxp_functions_0_aadd_17_a152;
wire fxp_functions_0_aadd_17_a156_sumout;
wire fxp_functions_0_aadd_17_a162_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq;
wire fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aadd_13_a1_sumout;
wire fxp_functions_0_aadd_13_a2;
wire fxp_functions_0_aadd_13_a6_sumout;
wire fxp_functions_0_aadd_13_a7;
wire fxp_functions_0_aadd_13_a11_sumout;
wire fxp_functions_0_aadd_13_a12;
wire fxp_functions_0_aadd_13_a16_sumout;
wire fxp_functions_0_aadd_13_a17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aadd_13_a21_sumout;
wire fxp_functions_0_aadd_13_a22;
wire fxp_functions_0_aadd_13_a26_sumout;
wire fxp_functions_0_aadd_13_a27;
wire fxp_functions_0_aadd_13_a31_sumout;
wire fxp_functions_0_aadd_13_a32;
wire fxp_functions_0_aadd_13_a36_sumout;
wire fxp_functions_0_aadd_13_a37;
wire fxp_functions_0_aadd_13_a41_sumout;
wire fxp_functions_0_aadd_13_a42;
wire fxp_functions_0_aadd_13_a46_sumout;
wire fxp_functions_0_aadd_13_a47;
wire fxp_functions_0_aadd_13_a51_sumout;
wire fxp_functions_0_aadd_13_a52;
wire fxp_functions_0_aadd_13_a56_sumout;
wire fxp_functions_0_aadd_13_a57;
wire fxp_functions_0_aadd_13_a61_sumout;
wire fxp_functions_0_aadd_13_a62;
wire fxp_functions_0_aadd_13_a66_sumout;
wire fxp_functions_0_aadd_13_a67;
wire fxp_functions_0_aadd_13_a71_sumout;
wire fxp_functions_0_aadd_13_a72;
wire fxp_functions_0_aadd_13_a76_sumout;
wire fxp_functions_0_aadd_13_a77;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aadd_13_a81_sumout;
wire fxp_functions_0_aadd_13_a82;
wire fxp_functions_0_aadd_13_a86_sumout;
wire fxp_functions_0_aadd_13_a87;
wire fxp_functions_0_aadd_13_a91_sumout;
wire fxp_functions_0_aadd_13_a92;
wire fxp_functions_0_aadd_13_a96_sumout;
wire fxp_functions_0_aadd_13_a97;
wire fxp_functions_0_aadd_13_a101_sumout;
wire fxp_functions_0_aadd_13_a102;
wire fxp_functions_0_aadd_13_a106_sumout;
wire fxp_functions_0_aadd_13_a107;
wire fxp_functions_0_aadd_13_a111_sumout;
wire fxp_functions_0_aadd_13_a112;
wire fxp_functions_0_aadd_13_a116_sumout;
wire fxp_functions_0_aadd_13_a117;
wire fxp_functions_0_aadd_13_a121_sumout;
wire fxp_functions_0_aadd_13_a122;
wire fxp_functions_0_aadd_13_a126_sumout;
wire fxp_functions_0_aadd_13_a127;
wire fxp_functions_0_aadd_13_a131_sumout;
wire fxp_functions_0_aadd_13_a132;
wire fxp_functions_0_aadd_13_a136_sumout;
wire fxp_functions_0_aadd_13_a137;
wire fxp_functions_0_aadd_13_a141_sumout;
wire fxp_functions_0_aadd_13_a142;
wire fxp_functions_0_aadd_13_a146_sumout;
wire fxp_functions_0_aadd_13_a147;
wire fxp_functions_0_aadd_13_a151_sumout;
wire fxp_functions_0_aadd_13_a152;
wire fxp_functions_0_aadd_13_a156_sumout;
wire fxp_functions_0_aadd_13_a157;
wire fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a_aq;
wire fxp_functions_0_aadd_13_a161_sumout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aadd_13_a166_sumout;
wire fxp_functions_0_aadd_13_a167;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a0_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a1_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a2_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a3_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a4_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a5_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a6_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a7_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a8_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a9_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a10_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a11_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a12_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a13_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a14_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a15_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a16_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a17_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a18_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a19_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a20_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a21_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a22_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a23_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a24_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a25_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a26_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a27_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a28_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a29_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a30_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA31;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA32;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA33;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA34;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA35;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a0_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a1_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a2_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a3_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a4_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a5_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a6_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a7_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a8_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a9_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a10_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a11_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a12_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a13_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a14_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a15_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a16_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a17_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a18_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a19_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a20_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a21_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a22_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a23_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a24_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a25_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a26_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a27_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a28_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a29_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a30_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a31_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a32_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a33_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA34;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA35;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a0_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a1_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a2_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a3_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a4_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a5_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a6_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a7_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a8_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a9_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a10_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a11_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a12_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a13_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a14_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a15_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a16_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a17_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a18_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a19_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a20_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a21_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a22_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a23_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a24_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a25_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a26_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a27_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a28_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a29_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a30_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a31_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a32_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a33_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a34_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a35_a;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_aadd_13_a172_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aadd_13_a177_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a_aq;
wire fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq;
wire fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq;
wire fxp_functions_0_aadd_13_a182_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq;
wire fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a_aq;
wire fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aadd_12_a1_sumout;
wire fxp_functions_0_aadd_12_a2;
wire fxp_functions_0_aadd_12_a6_sumout;
wire fxp_functions_0_aadd_12_a7;
wire fxp_functions_0_aadd_12_a11_sumout;
wire fxp_functions_0_aadd_12_a12;
wire fxp_functions_0_aadd_12_a16_sumout;
wire fxp_functions_0_aadd_12_a17;
wire fxp_functions_0_aadd_12_a21_sumout;
wire fxp_functions_0_aadd_12_a22;
wire fxp_functions_0_aadd_12_a26_sumout;
wire fxp_functions_0_aadd_12_a27;
wire fxp_functions_0_aadd_12_a31_sumout;
wire fxp_functions_0_aadd_12_a32;
wire fxp_functions_0_aadd_12_a36_sumout;
wire fxp_functions_0_aadd_12_a37;
wire fxp_functions_0_aadd_12_a41_sumout;
wire fxp_functions_0_aadd_12_a42;
wire fxp_functions_0_aadd_12_a46_sumout;
wire fxp_functions_0_aadd_12_a47;
wire fxp_functions_0_aadd_12_a51_sumout;
wire fxp_functions_0_aadd_12_a52;
wire fxp_functions_0_aadd_12_a56_sumout;
wire fxp_functions_0_aadd_12_a57;
wire fxp_functions_0_aadd_12_a61_sumout;
wire fxp_functions_0_aadd_12_a62;
wire fxp_functions_0_aadd_12_a66_sumout;
wire fxp_functions_0_aadd_12_a67;
wire fxp_functions_0_aadd_12_a71_sumout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq;
wire fxp_functions_0_aadd_12_a76_sumout;
wire fxp_functions_0_aadd_12_a77;
wire fxp_functions_0_aadd_12_a81_sumout;
wire fxp_functions_0_aadd_12_a82;
wire fxp_functions_0_aadd_12_a86_sumout;
wire fxp_functions_0_aadd_12_a87;
wire fxp_functions_0_aadd_12_a91_sumout;
wire fxp_functions_0_aadd_12_a92;
wire fxp_functions_0_aadd_12_a96_sumout;
wire fxp_functions_0_aadd_12_a97;
wire fxp_functions_0_aadd_12_a101_sumout;
wire fxp_functions_0_aadd_12_a102;
wire fxp_functions_0_aadd_12_a106_sumout;
wire fxp_functions_0_aadd_12_a107;
wire fxp_functions_0_aadd_12_a111_sumout;
wire fxp_functions_0_aadd_12_a112;
wire fxp_functions_0_aadd_12_a116_sumout;
wire fxp_functions_0_aadd_12_a117;
wire fxp_functions_0_aadd_12_a121_sumout;
wire fxp_functions_0_aadd_12_a122;
wire fxp_functions_0_aadd_12_a126_sumout;
wire fxp_functions_0_aadd_12_a127;
wire fxp_functions_0_aadd_12_a131_sumout;
wire fxp_functions_0_aadd_12_a132;
wire fxp_functions_0_aadd_12_a136_sumout;
wire fxp_functions_0_aadd_12_a137;
wire fxp_functions_0_aadd_12_a141_sumout;
wire fxp_functions_0_aadd_12_a142;
wire fxp_functions_0_aadd_12_a146_sumout;
wire fxp_functions_0_aadd_12_a147;
wire fxp_functions_0_aadd_12_a151_sumout;
wire fxp_functions_0_aadd_12_a152;
wire fxp_functions_0_aadd_12_a156_sumout;
wire fxp_functions_0_aadd_12_a157;
wire fxp_functions_0_aadd_12_a161_sumout;
wire fxp_functions_0_aadd_12_a162;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a_aq;
wire fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a_aq;
wire fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a_aq;
wire fxp_functions_0_aadd_13_a187_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a_aq;
wire fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a_aq;
wire fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a24_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a25_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a26_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a27_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a28_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a29_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a30_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a31_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT19;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a_aq;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a30_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a31_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a32_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a33_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a34_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a35_a;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a36_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fxp_functions_0_aadd_12_a167_cout;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a_aq;
wire fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a_aq;
wire fxp_functions_0_aadd_13_a192_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a_aq;
wire fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a_aq;
wire fxp_functions_0_aadd_9_a1_sumout;
wire fxp_functions_0_aadd_9_a2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aadd_9_a6_sumout;
wire fxp_functions_0_aadd_9_a7;
wire fxp_functions_0_aadd_9_a11_sumout;
wire fxp_functions_0_aadd_9_a12;
wire fxp_functions_0_aadd_9_a16_sumout;
wire fxp_functions_0_aadd_9_a17;
wire fxp_functions_0_aadd_9_a21_sumout;
wire fxp_functions_0_aadd_9_a22;
wire fxp_functions_0_aadd_9_a26_sumout;
wire fxp_functions_0_aadd_9_a27;
wire fxp_functions_0_aadd_9_a31_sumout;
wire fxp_functions_0_aadd_9_a32;
wire fxp_functions_0_aadd_9_a36_sumout;
wire fxp_functions_0_aadd_9_a41_sumout;
wire fxp_functions_0_aadd_9_a42;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fxp_functions_0_aadd_12_a172_cout;
wire fxp_functions_0_aadd_9_a46_sumout;
wire fxp_functions_0_aadd_9_a47;
wire fxp_functions_0_aadd_9_a51_sumout;
wire fxp_functions_0_aadd_9_a52;
wire fxp_functions_0_aadd_9_a56_sumout;
wire fxp_functions_0_aadd_9_a57;
wire fxp_functions_0_aadd_9_a61_sumout;
wire fxp_functions_0_aadd_9_a62;
wire fxp_functions_0_aadd_9_a66_sumout;
wire fxp_functions_0_aadd_9_a67;
wire fxp_functions_0_aadd_9_a71_sumout;
wire fxp_functions_0_aadd_9_a72;
wire fxp_functions_0_aadd_9_a76_sumout;
wire fxp_functions_0_aadd_9_a77;
wire fxp_functions_0_aadd_9_a81_sumout;
wire fxp_functions_0_aadd_9_a82;
wire fxp_functions_0_aadd_9_a86_sumout;
wire fxp_functions_0_aadd_9_a87;
wire fxp_functions_0_aadd_9_a91_sumout;
wire fxp_functions_0_aadd_9_a92;
wire fxp_functions_0_aadd_9_a96_sumout;
wire fxp_functions_0_aadd_9_a97;
wire fxp_functions_0_aadd_9_a101_sumout;
wire fxp_functions_0_aadd_9_a102;
wire fxp_functions_0_aadd_9_a106_sumout;
wire fxp_functions_0_aadd_9_a107;
wire fxp_functions_0_aadd_9_a111_sumout;
wire fxp_functions_0_aadd_9_a112;
wire fxp_functions_0_aadd_9_a116_sumout;
wire fxp_functions_0_aadd_9_a117;
wire fxp_functions_0_aadd_9_a121_sumout;
wire fxp_functions_0_aadd_9_a122;
wire fxp_functions_0_aadd_9_a126_sumout;
wire fxp_functions_0_aadd_9_a127;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a_aq;
wire fxp_functions_0_aadd_13_a197_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a_aq;
wire fxp_functions_0_aadd_9_a131_sumout;
wire fxp_functions_0_aadd_9_a132;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fxp_functions_0_aadd_12_a177_cout;
wire fxp_functions_0_aadd_13_a202_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a0_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a1_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a2_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a3_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a4_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a5_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a6_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a7_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a8_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a9_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a10_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a11_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a12_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a13_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a14_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a15_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a16_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a17_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a18_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a19_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a20_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a21_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a22_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a23_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a24_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a25_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a26_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a27_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a28_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a29_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a30_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a31_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a32_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a33_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a34_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a35_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a36_a;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a0_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a1_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a2_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a3_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a4_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a5_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a6_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a7_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a8_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a9_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a10_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a11_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a12_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a13_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a14_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a15_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a16_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a17_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a18_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a19_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a20_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a21_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a22_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a23_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a24_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a25_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a26_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a27_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a28_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a29_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a30_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a31_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a32_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a33_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a34_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a35_a;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fxp_functions_0_aadd_9_a136_sumout;
wire fxp_functions_0_aadd_9_a137;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fxp_functions_0_aadd_12_a182_cout;
wire fxp_functions_0_aadd_13_a207_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aadd_9_a141_sumout;
wire fxp_functions_0_aadd_9_a142;
wire fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a_aq;
wire fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fxp_functions_0_aadd_13_a212_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a_aq;
wire fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a_aq;
wire fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a_aq;
wire fxp_functions_0_aadd_9_a146_sumout;
wire fxp_functions_0_aadd_9_a147;
wire fxp_functions_0_aadd_13_a217_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq;
wire fxp_functions_0_aadd_8_a1_sumout;
wire fxp_functions_0_aadd_8_a2;
wire fxp_functions_0_aadd_8_a6_sumout;
wire fxp_functions_0_aadd_8_a7;
wire fxp_functions_0_aadd_8_a11_sumout;
wire fxp_functions_0_aadd_8_a12;
wire fxp_functions_0_aadd_8_a16_sumout;
wire fxp_functions_0_aadd_8_a17;
wire fxp_functions_0_aadd_8_a21_sumout;
wire fxp_functions_0_aadd_8_a22;
wire fxp_functions_0_aadd_8_a26_sumout;
wire fxp_functions_0_aadd_8_a27;
wire fxp_functions_0_aadd_8_a31_sumout;
wire fxp_functions_0_aadd_8_a32;
wire fxp_functions_0_aadd_8_a36_sumout;
wire fxp_functions_0_aadd_8_a37;
wire fxp_functions_0_aadd_8_a41_sumout;
wire fxp_functions_0_aadd_8_a42;
wire fxp_functions_0_aadd_8_a46_sumout;
wire fxp_functions_0_aadd_8_a47;
wire fxp_functions_0_aadd_8_a51_sumout;
wire fxp_functions_0_aadd_8_a52;
wire fxp_functions_0_aadd_8_a56_sumout;
wire fxp_functions_0_aadd_8_a57;
wire fxp_functions_0_aadd_8_a61_sumout;
wire fxp_functions_0_aadd_8_a62;
wire fxp_functions_0_aadd_8_a66_sumout;
wire fxp_functions_0_aadd_8_a67;
wire fxp_functions_0_aadd_8_a71_sumout;
wire fxp_functions_0_aadd_8_a72;
wire fxp_functions_0_aadd_8_a76_sumout;
wire fxp_functions_0_aadd_8_a77;
wire fxp_functions_0_aadd_8_a81_sumout;
wire fxp_functions_0_aadd_8_a82;
wire fxp_functions_0_aadd_8_a86_sumout;
wire fxp_functions_0_aadd_8_a87;
wire fxp_functions_0_aadd_8_a91_sumout;
wire fxp_functions_0_aadd_8_a92;
wire fxp_functions_0_aadd_8_a96_sumout;
wire fxp_functions_0_aadd_8_a97;
wire fxp_functions_0_aadd_8_a101_sumout;
wire fxp_functions_0_aadd_8_a102;
wire fxp_functions_0_aadd_8_a106_sumout;
wire fxp_functions_0_aadd_8_a107;
wire fxp_functions_0_aadd_8_a111_sumout;
wire fxp_functions_0_aadd_8_a112;
wire fxp_functions_0_aadd_8_a116_sumout;
wire fxp_functions_0_aadd_8_a117;
wire fxp_functions_0_aadd_8_a121_sumout;
wire fxp_functions_0_aadd_8_a122;
wire fxp_functions_0_aadd_8_a126_sumout;
wire fxp_functions_0_aadd_8_a127;
wire fxp_functions_0_aadd_8_a131_sumout;
wire fxp_functions_0_aadd_8_a132;
wire fxp_functions_0_aadd_8_a136_sumout;
wire fxp_functions_0_aadd_8_a137;
wire fxp_functions_0_aadd_8_a141_sumout;
wire fxp_functions_0_aadd_8_a142;
wire fxp_functions_0_aadd_8_a146_sumout;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aadd_9_a152_cout;
wire fxp_functions_0_aadd_13_a222_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a0_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a1_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a2_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a3_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a4_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a5_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a6_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a7_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a8_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a9_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a10_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a11_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a12_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a13_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a14_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a15_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a16_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a17_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a18_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a19_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a20_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a21_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a22_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a23_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a24_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a25_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a26_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a27_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a28_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a29_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a30_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a31_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a32_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a33_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a34_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a35_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a36_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a37_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a38_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a39_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a40_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a41_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a42_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a43_a;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a;
wire fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a_aq;
wire fxp_functions_0_aadd_9_a157_cout;
wire fxp_functions_0_aadd_13_a227_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a_aq;
wire fxp_functions_0_aadd_9_a162_cout;
wire fxp_functions_0_aadd_13_a232_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a_aq;
wire fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a_aq;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a_aq;
wire fxp_functions_0_aadd_9_a167_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a_aq;
wire fxp_functions_0_aadd_7_a1_sumout;
wire fxp_functions_0_aadd_7_a2;
wire fxp_functions_0_aadd_7_a6_sumout;
wire fxp_functions_0_aadd_7_a7;
wire fxp_functions_0_aadd_7_a11_sumout;
wire fxp_functions_0_aadd_7_a12;
wire fxp_functions_0_aadd_7_a16_sumout;
wire fxp_functions_0_aadd_7_a17;
wire fxp_functions_0_aadd_7_a21_sumout;
wire fxp_functions_0_aadd_7_a22;
wire fxp_functions_0_aadd_7_a26_sumout;
wire fxp_functions_0_aadd_7_a27;
wire fxp_functions_0_aadd_7_a31_sumout;
wire fxp_functions_0_aadd_7_a32;
wire fxp_functions_0_aadd_7_a36_sumout;
wire fxp_functions_0_aadd_7_a37;
wire fxp_functions_0_aadd_7_a41_sumout;
wire fxp_functions_0_aadd_7_a42;
wire fxp_functions_0_aadd_7_a46_sumout;
wire fxp_functions_0_aadd_7_a47;
wire fxp_functions_0_aadd_7_a51_sumout;
wire fxp_functions_0_aadd_7_a52;
wire fxp_functions_0_aadd_7_a56_sumout;
wire fxp_functions_0_aadd_7_a57;
wire fxp_functions_0_aadd_7_a61_sumout;
wire fxp_functions_0_aadd_7_a62;
wire fxp_functions_0_aadd_7_a66_sumout;
wire fxp_functions_0_aadd_7_a67;
wire fxp_functions_0_aadd_7_a71_sumout;
wire fxp_functions_0_aadd_7_a72;
wire fxp_functions_0_aadd_7_a76_sumout;
wire fxp_functions_0_aadd_7_a77;
wire fxp_functions_0_aadd_7_a81_sumout;
wire fxp_functions_0_aadd_7_a82;
wire fxp_functions_0_aadd_7_a86_sumout;
wire fxp_functions_0_aadd_7_a87;
wire fxp_functions_0_aadd_7_a91_sumout;
wire fxp_functions_0_aadd_7_a92;
wire fxp_functions_0_aadd_7_a96_sumout;
wire fxp_functions_0_aadd_7_a97;
wire fxp_functions_0_aadd_7_a101_sumout;
wire fxp_functions_0_aadd_7_a102;
wire fxp_functions_0_aadd_7_a106_sumout;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a_aq;
wire fxp_functions_0_aadd_9_a172_cout;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a0_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a1_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a2_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a3_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a4_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a5_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a6_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a7_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a8_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a9_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a10_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a11_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a12_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a13_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a14_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a15_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a16_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a17_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a18_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a19_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a20_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a21_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a22_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a23_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a24_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a25_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a26_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a27_a;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA28;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA29;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA30;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA31;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA32;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA33;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA34;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA35;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA36;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA37;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA38;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA39;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA40;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA41;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA42;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA43;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA44;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA45;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA46;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA47;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA48;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA49;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA50;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA51;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA52;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA53;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA54;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA55;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA56;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA57;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA58;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA59;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA60;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA61;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA62;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA63;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a;
wire fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a_aq;
wire fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a_aq;
wire fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a_aq;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a;
wire fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a_aq;
wire fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a_aq;
wire fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a_aq;
wire fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a_aq;
wire fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a_aq;
wire fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a_aq;
wire fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a_aq;
wire fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a_aq;
wire fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a_aq;
wire fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a_aq;
wire fxp_functions_0_aMux_99_a2_cout;
wire fxp_functions_0_aMux_99_a6_sumout;
wire fxp_functions_0_aMux_99_a7;
wire fxp_functions_0_aMux_100_a1_sumout;
wire fxp_functions_0_aMux_100_a2;
wire fxp_functions_0_aMux_101_a1_sumout;
wire fxp_functions_0_aMux_101_a2;
wire fxp_functions_0_aMux_102_a1_sumout;
wire fxp_functions_0_aMux_102_a2;
wire fxp_functions_0_aMux_103_a1_sumout;
wire fxp_functions_0_aMux_103_a2;
wire fxp_functions_0_aMux_104_a1_sumout;
wire fxp_functions_0_aMux_104_a2;
wire fxp_functions_0_aMux_105_a1_sumout;
wire fxp_functions_0_aMux_105_a2;
wire fxp_functions_0_aMux_106_a1_sumout;
wire fxp_functions_0_aMux_106_a2;
wire fxp_functions_0_aMux_107_a1_sumout;
wire fxp_functions_0_aMux_107_a2;
wire fxp_functions_0_aMux_108_a1_sumout;
wire fxp_functions_0_aMux_108_a2;
wire fxp_functions_0_aMux_109_a1_sumout;
wire fxp_functions_0_aMux_109_a2;
wire fxp_functions_0_aMux_110_a1_sumout;
wire fxp_functions_0_aMux_110_a2;
wire fxp_functions_0_aMux_111_a1_sumout;
wire fxp_functions_0_aMux_111_a2;
wire fxp_functions_0_aMux_112_a1_sumout;
wire fxp_functions_0_aMux_112_a2;
wire fxp_functions_0_aMux_113_a1_sumout;
wire fxp_functions_0_aMux_113_a2;
wire fxp_functions_0_aMux_114_a1_sumout;
wire fxp_functions_0_aMux_114_a2;
wire fxp_functions_0_aMux_115_a1_sumout;
wire fxp_functions_0_aMux_115_a2;
wire fxp_functions_0_aMux_116_a1_sumout;
wire fxp_functions_0_aMux_116_a2;
wire fxp_functions_0_aMux_117_a1_sumout;
wire fxp_functions_0_aMux_118_a2_cout;
wire fxp_functions_0_aMux_118_a6_sumout;
wire fxp_functions_0_aMux_118_a7;
wire fxp_functions_0_aMux_119_a1_sumout;
wire fxp_functions_0_aMux_119_a2;
wire fxp_functions_0_aMux_120_a1_sumout;
wire fxp_functions_0_aMux_120_a2;
wire fxp_functions_0_aMux_121_a1_sumout;
wire fxp_functions_0_aMux_121_a2;
wire fxp_functions_0_aMux_122_a1_sumout;
wire fxp_functions_0_aMux_122_a2;
wire fxp_functions_0_aMux_123_a1_sumout;
wire fxp_functions_0_aMux_123_a2;
wire fxp_functions_0_aMux_124_a1_sumout;
wire fxp_functions_0_aMux_124_a2;
wire fxp_functions_0_aMux_125_a1_sumout;
wire fxp_functions_0_aMux_125_a2;
wire fxp_functions_0_ai8489_a13_sumout;
wire fxp_functions_0_ai8489_a14;
wire fxp_functions_0_ai8489_a18_sumout;
wire fxp_functions_0_ai8489_a19;
wire fxp_functions_0_ai8489_a23_sumout;
wire fxp_functions_0_ai8489_a24;
wire fxp_functions_0_ai8489_a28_sumout;
wire fxp_functions_0_aMux_48_a2_cout;
wire fxp_functions_0_aMux_48_a6_sumout;
wire fxp_functions_0_aMux_48_a7;
wire fxp_functions_0_aMux_44_a1_sumout;
wire fxp_functions_0_aMux_44_a2;
wire fxp_functions_0_aMux_40_a19_sumout;
wire fxp_functions_0_aMux_50_a2_cout;
wire fxp_functions_0_aMux_50_a6_sumout;
wire fxp_functions_0_aMux_50_a7;
wire fxp_functions_0_aMux_46_a1_sumout;
wire fxp_functions_0_aMux_46_a2;
wire fxp_functions_0_aMux_42_a1_sumout;
wire fxp_functions_0_aMux_49_a2_cout;
wire fxp_functions_0_aMux_49_a6_sumout;
wire fxp_functions_0_aMux_49_a7;
wire fxp_functions_0_aMux_45_a1_sumout;
wire fxp_functions_0_aMux_45_a2;
wire fxp_functions_0_aMux_41_a1_sumout;
wire fxp_functions_0_aMux_51_a2_cout;
wire fxp_functions_0_aMux_51_a6_sumout;
wire fxp_functions_0_aMux_51_a7;
wire fxp_functions_0_aMux_47_a1_sumout;
wire fxp_functions_0_aMux_47_a2;
wire fxp_functions_0_aMux_43_a1_sumout;
wire fxp_functions_0_ai6615_a2_cout;
wire fxp_functions_0_ai6615_a6_sumout;
wire fxp_functions_0_ai6615_a7;
wire fxp_functions_0_ai6615_a11_sumout;
wire fxp_functions_0_ai6615_a12;
wire fxp_functions_0_ai6615_a16_sumout;
wire fxp_functions_0_ai6615_a17;
wire fxp_functions_0_ai6615_a21_sumout;
wire fxp_functions_0_ai6615_a22;
wire fxp_functions_0_ai6615_a26_sumout;
wire fxp_functions_0_ai6615_a27;
wire fxp_functions_0_ai6615_a31_sumout;
wire fxp_functions_0_ai6615_a32;
wire fxp_functions_0_ai6615_a36_sumout;
wire fxp_functions_0_ai6615_a37;
wire fxp_functions_0_ai6615_a41_sumout;
wire fxp_functions_0_ai6615_a42;
wire fxp_functions_0_ai6615_a46_sumout;
wire fxp_functions_0_ai6615_a47;
wire fxp_functions_0_ai6615_a51_sumout;
wire fxp_functions_0_ai6615_a52;
wire fxp_functions_0_ai6615_a56_sumout;
wire fxp_functions_0_ai6615_a57;
wire fxp_functions_0_ai6615_a61_sumout;
wire fxp_functions_0_ai6615_a62;
wire fxp_functions_0_ai6615_a66_sumout;
wire fxp_functions_0_ai6615_a67;
wire fxp_functions_0_ai6615_a71_sumout;
wire fxp_functions_0_ai6615_a72;
wire fxp_functions_0_ai6615_a76_sumout;
wire fxp_functions_0_ai6615_a77;
wire fxp_functions_0_ai6615_a81_sumout;
wire fxp_functions_0_ai6615_a82;
wire fxp_functions_0_ai6615_a86_sumout;
wire fxp_functions_0_ai6615_a87;
wire fxp_functions_0_ai6615_a91_sumout;
wire fxp_functions_0_ai6615_a92;
wire fxp_functions_0_ai6615_a96_sumout;
wire fxp_functions_0_ai6615_a102_cout;
wire fxp_functions_0_ai6615_a106_sumout;
wire fxp_functions_0_ai6615_a107;
wire fxp_functions_0_aMux_72_a2_sumout;
wire fxp_functions_0_aMux_72_a3;
wire fxp_functions_0_aMux_72_a7_sumout;
wire fxp_functions_0_aMux_72_a8;
wire fxp_functions_0_aMux_72_a12_sumout;
wire fxp_functions_0_aMux_72_a13;
wire fxp_functions_0_aMux_72_a17_sumout;
wire fxp_functions_0_aMux_72_a18;
wire fxp_functions_0_aMux_72_a22_sumout;
wire fxp_functions_0_aMux_72_a23;
wire fxp_functions_0_aMux_72_a27_sumout;
wire fxp_functions_0_aMux_72_a28;
wire fxp_functions_0_aMux_72_a32_sumout;
wire fxp_functions_0_aMux_64_a1_combout;
wire fxp_functions_0_aMux_32_a3_combout;
wire fxp_functions_0_aMux_64_a6_combout;
wire fxp_functions_0_aMux_40_a23_combout;
wire fxp_functions_0_ai8489_a34_combout;
wire fxp_functions_0_ai8489_a39_combout;
wire fxp_functions_0_ai8489_a44_combout;
wire fxp_functions_0_ai8489_a49_combout;
wire fxp_functions_0_ai8489_a54_combout;
wire fxp_functions_0_ai8489_a59_combout;
wire fxp_functions_0_ai8489_a64_combout;
wire fxp_functions_0_ai8489_a69_combout;
wire fxp_functions_0_ai8489_a74_combout;
wire fxp_functions_0_ai8489_a79_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30_combout;
wire fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31_combout;
wire fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a_aq;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a_aq;
wire fxp_functions_0_aMux_177_a0_combout;
wire fxp_functions_0_ai8489_a0_combout;
wire fxp_functions_0_ai8489_a1_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a_aq;
wire fxp_functions_0_areduce_nor_0_a0_combout;
wire fxp_functions_0_areduce_nor_0_a1_combout;
wire fxp_functions_0_areduce_nor_0_a2_combout;
wire fxp_functions_0_areduce_nor_0_a3_combout;
wire fxp_functions_0_areduce_nor_0_a4_combout;
wire fxp_functions_0_areduce_nor_0_a5_combout;
wire fxp_functions_0_areduce_nor_0_acombout;
wire fxp_functions_0_aMux_176_a0_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1_combout;
wire fxp_functions_0_ai8489_a2_combout;
wire fxp_functions_0_ai8489_a3_combout;
wire fxp_functions_0_ai8489_a4_combout;
wire fxp_functions_0_aMux_98_a0_combout;
wire fxp_functions_0_aMux_175_a0_combout;
wire fxp_functions_0_ai8489_a5_combout;
wire fxp_functions_0_aMux_97_a1_combout;
wire fxp_functions_0_aMux_174_a0_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout;
wire fxp_functions_0_aMux_96_a0_combout;
wire fxp_functions_0_aMux_173_a0_combout;
wire fxp_functions_0_aMux_172_a0_combout;
wire fxp_functions_0_aMux_171_a0_combout;
wire fxp_functions_0_aMux_170_a0_combout;
wire fxp_functions_0_aMux_169_a0_combout;
wire fxp_functions_0_aMux_168_a1_combout;
wire fxp_functions_0_aMux_167_a1_combout;
wire fxp_functions_0_aMux_166_a1_combout;
wire fxp_functions_0_ai8489_a6_combout;
wire fxp_functions_0_aMux_165_a1_combout;
wire fxp_functions_0_ai8489_a7_combout;
wire fxp_functions_0_aMux_162_a0_combout;
wire fxp_functions_0_aMux_164_a0_combout;
wire fxp_functions_0_aMux_163_a0_combout;
wire fxp_functions_0_aMux_178_a0_combout;
wire fxp_functions_0_aMux_162_a1_combout;
wire fxp_functions_0_ai8489_a8_combout;
wire fxp_functions_0_ai8489_a9_combout;
wire fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout;
wire fxp_functions_0_ai8489_a10_combout;
wire fxp_functions_0_ai8489_a11_combout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq;
wire fxp_functions_0_ai8103_a0_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1_combout;
wire fxp_functions_0_ai8150_a0_combout;
wire fxp_functions_0_ai8150_a1_combout;
wire fxp_functions_0_ai8150_a2_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4_combout;
wire fxp_functions_0_areduce_nor_21_acombout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_ai8126_a0_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0_combout;
wire fxp_functions_0_aadd_15_a0_combout;
wire fxp_functions_0_ai8126_a1_combout;
wire fxp_functions_0_ai8126_a2_combout;
wire fxp_functions_0_ai8126_a3_combout;
wire fxp_functions_0_ai6816_a0_combout;
wire fxp_functions_0_ai6816_a1_combout;
wire fxp_functions_0_ai6816_a2_combout;
wire fxp_functions_0_ai6816_a3_combout;
wire fxp_functions_0_ai6816_a4_combout;
wire fxp_functions_0_ai6816_a5_combout;
wire fxp_functions_0_ai6816_a6_combout;
wire fxp_functions_0_ai6816_a7_combout;
wire fxp_functions_0_ai6816_a8_combout;
wire fxp_functions_0_ai6816_a9_combout;
wire fxp_functions_0_ai6816_a10_combout;
wire fxp_functions_0_ai6816_a11_combout;
wire fxp_functions_0_ai6816_a12_combout;
wire fxp_functions_0_ai6816_a13_combout;
wire fxp_functions_0_ai6816_a14_combout;
wire fxp_functions_0_ai6816_a15_combout;
wire fxp_functions_0_ai6816_a16_combout;
wire fxp_functions_0_ai6816_a17_combout;
wire fxp_functions_0_ai6816_a18_combout;
wire fxp_functions_0_ai6816_a19_combout;
wire fxp_functions_0_ai6816_a20_combout;
wire fxp_functions_0_ai6816_a21_combout;
wire fxp_functions_0_ai6816_a22_combout;
wire fxp_functions_0_ai6816_a23_combout;
wire fxp_functions_0_ai6816_a24_combout;
wire fxp_functions_0_ai6816_a25_combout;
wire fxp_functions_0_ai6816_a26_combout;
wire fxp_functions_0_ai6816_a27_combout;
wire fxp_functions_0_ai6816_a28_combout;
wire fxp_functions_0_ai6816_a29_combout;
wire fxp_functions_0_ai6816_a30_combout;
wire fxp_functions_0_ai6816_a31_combout;
wire fxp_functions_0_ai6816_a32_combout;
wire fxp_functions_0_areduce_nor_10_a1_combout;
wire fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0_combout;
wire fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1_combout;
wire fxp_functions_0_areduce_nor_9_acombout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_areduce_nor_17_acombout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_ai3244_a1_combout;
wire fxp_functions_0_ai3244_a2_combout;
wire fxp_functions_0_ai3244_a3_combout;
wire fxp_functions_0_ai3244_a4_combout;
wire fxp_functions_0_ai3244_a5_combout;
wire fxp_functions_0_ai3244_a6_combout;
wire fxp_functions_0_ai3244_a7_combout;
wire fxp_functions_0_ai3244_a8_combout;
wire fxp_functions_0_ai3244_a9_combout;
wire fxp_functions_0_ai3244_a10_combout;
wire fxp_functions_0_ai3244_a11_combout;
wire fxp_functions_0_ai3244_a12_combout;
wire fxp_functions_0_areduce_nor_8_acombout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_areduce_nor_7_a0_combout;
wire fxp_functions_0_areduce_nor_7_a1_combout;
wire fxp_functions_0_areduce_nor_7_a2_combout;
wire fxp_functions_0_areduce_nor_7_a3_combout;
wire fxp_functions_0_areduce_nor_7_a4_combout;
wire fxp_functions_0_areduce_nor_7_a5_combout;
wire fxp_functions_0_areduce_nor_7_acombout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq;
wire fxp_functions_0_ai1590_a0_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq;
wire fxp_functions_0_ai3159_a1_combout;
wire fxp_functions_0_ai3159_a2_combout;
wire fxp_functions_0_ai3159_a3_combout;
wire fxp_functions_0_ai3159_a4_combout;
wire fxp_functions_0_ai3159_a5_combout;
wire fxp_functions_0_ai3159_a6_combout;
wire fxp_functions_0_ai3159_a7_combout;
wire fxp_functions_0_ai3159_a8_combout;
wire fxp_functions_0_ai3159_a9_combout;
wire fxp_functions_0_ai3159_a10_combout;
wire fxp_functions_0_ai3159_a11_combout;
wire fxp_functions_0_ai3159_a12_combout;
wire fxp_functions_0_ai3159_a13_combout;
wire fxp_functions_0_ai3159_a14_combout;
wire fxp_functions_0_ai3159_a15_combout;
wire fxp_functions_0_ai3159_a16_combout;
wire fxp_functions_0_ai3159_a17_combout;
wire fxp_functions_0_ai3159_a18_combout;
wire fxp_functions_0_ai3159_a19_combout;
wire fxp_functions_0_ai3159_a20_combout;
wire fxp_functions_0_ai3159_a21_combout;
wire fxp_functions_0_ai3159_a22_combout;
wire fxp_functions_0_ai3159_a23_combout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_areduce_nor_6_a0_combout;
wire fxp_functions_0_areduce_nor_6_a1_combout;
wire fxp_functions_0_areduce_nor_6_a2_combout;
wire fxp_functions_0_areduce_nor_6_a3_combout;
wire fxp_functions_0_areduce_nor_6_a4_combout;
wire fxp_functions_0_areduce_nor_6_a5_combout;
wire fxp_functions_0_areduce_nor_6_acombout;
wire fxp_functions_0_ai1731_a0_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1_combout;
wire fxp_functions_0_ai1731_a1_combout;
wire fxp_functions_0_ai1731_a2_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4_combout;
wire fxp_functions_0_areduce_nor_19_acombout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_aadd_0_a0_combout;
wire fxp_functions_0_aadd_0_a1_combout;
wire fxp_functions_0_aadd_0_a2_combout;
wire fxp_functions_0_aadd_0_a3_combout;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_areduce_nor_2_acombout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fxp_functions_0_ai6102_a0_combout;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0_combout;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1_combout;
wire fxp_functions_0_ai6157_a0_combout;
wire fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2_combout;
wire fxp_functions_0_areduce_nor_13_acombout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_ai6114_a0_combout;
wire fxp_functions_0_ai6114_a1_combout;
wire fxp_functions_0_ai6114_a2_combout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq;
wire fxp_functions_0_areduce_nor_14_acombout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_ai1992_a0_combout;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_ai3830_a0_combout;
wire fxp_functions_0_ai3830_a1_combout;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0_combout;
wire fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1_combout;
wire fxp_functions_0_areduce_nor_20_acombout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_ai1997_a0_combout;
wire fxp_functions_0_aadd_2_a0_combout;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a_aq;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a_aq;
wire fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fxp_functions_0_ai2020_a0_combout;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0_combout;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1_combout;
wire fxp_functions_0_ai3634_a0_combout;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2_combout;
wire fxp_functions_0_areduce_nor_4_acombout;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout;
wire fxp_functions_0_ai2032_a0_combout;
wire fxp_functions_0_ai2032_a1_combout;
wire fxp_functions_0_ai2032_a2_combout;
wire fxp_functions_0_aMux_8_a1_combout;
wire fxp_functions_0_aMux_16_a0_combout;
wire fxp_functions_0_aMux_12_a1_combout;
wire fxp_functions_0_aMux_20_a0_combout;
wire fxp_functions_0_aMux_10_a1_combout;
wire fxp_functions_0_aMux_18_a0_combout;
wire fxp_functions_0_aMux_14_a1_combout;
wire fxp_functions_0_aMux_22_a0_combout;
wire fxp_functions_0_aMux_9_a1_combout;
wire fxp_functions_0_aMux_17_a0_combout;
wire fxp_functions_0_aMux_13_a1_combout;
wire fxp_functions_0_aMux_21_a0_combout;
wire fxp_functions_0_aMux_11_a1_combout;
wire fxp_functions_0_aMux_19_a0_combout;
wire fxp_functions_0_aMux_15_a1_combout;
wire fxp_functions_0_aMux_23_a0_combout;
wire fxp_functions_0_aMux_40_a0_combout;
wire fxp_functions_0_aMux_40_a1_combout;
wire fxp_functions_0_aMux_40_a2_combout;
wire fxp_functions_0_aMux_40_a3_combout;
wire fxp_functions_0_aMux_40_a4_combout;
wire fxp_functions_0_aMux_40_a5_combout;
wire fxp_functions_0_aMux_40_a6_combout;
wire fxp_functions_0_aMux_40_a7_combout;
wire fxp_functions_0_aMux_40_a8_combout;
wire fxp_functions_0_aMux_32_a0_combout;
wire fxp_functions_0_aMux_32_a1_combout;
wire fxp_functions_0_aMux_40_a9_combout;
wire fxp_functions_0_aMux_40_a10_combout;
wire fxp_functions_0_aMux_40_a11_combout;
wire fxp_functions_0_aMux_40_a12_combout;
wire fxp_functions_0_aMux_40_a13_combout;
wire fxp_functions_0_aMux_40_a14_combout;
wire fxp_functions_0_aMux_40_a15_combout;
wire fxp_functions_0_aMux_40_a16_combout;
wire fxp_functions_0_aMux_72_a0_combout;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq;
wire fxp_functions_0_ai4258_a0_combout;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq;
wire fxp_functions_0_areduce_nor_5_acombout;
wire fxp_functions_0_aMux_30_a0_combout;
wire fxp_functions_0_aMux_26_a0_combout;
wire fxp_functions_0_aMux_54_a0_combout;
wire fxp_functions_0_aMux_94_a1_combout;
wire fxp_functions_0_aMux_56_a1_combout;
wire fxp_functions_0_aMux_31_a0_combout;
wire fxp_functions_0_aMux_27_a0_combout;
wire fxp_functions_0_aMux_55_a0_combout;
wire fxp_functions_0_aMux_57_a1_combout;
wire fxp_functions_0_aMux_29_a0_combout;
wire fxp_functions_0_aMux_25_a0_combout;
wire fxp_functions_0_aMux_53_a0_combout;
wire fxp_functions_0_aMux_28_a0_combout;
wire fxp_functions_0_aMux_24_a0_combout;
wire fxp_functions_0_aMux_52_a0_combout;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0_combout;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1_combout;
wire fxp_functions_0_ai4289_a0_combout;
wire fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2_combout;
wire fxp_functions_0_areduce_nor_11_acombout;
wire fxp_functions_0_aMux_63_a0_combout;
wire fxp_functions_0_aMux_61_a0_combout;
wire fxp_functions_0_aMux_62_a0_combout;
wire fxp_functions_0_aMux_93_a0_combout;
wire fxp_functions_0_aMux_60_a0_combout;
wire fxp_functions_0_aMux_59_a1_combout;
wire fxp_functions_0_aMux_58_a1_combout;
wire fxp_functions_0_ai4270_a0_combout;
wire fxp_functions_0_ai4270_a1_combout;
wire fxp_functions_0_ai4270_a2_combout;
wire fxp_functions_0_aMux_95_a0_combout;
wire fxp_functions_0_aMux_94_a2_combout;
wire fxp_functions_0_areduce_nor_12_acombout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7_combout;
wire fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0_combout;
wire fxp_functions_0_aMux_32_a2_combout;
wire fxp_functions_0_aMux_40_a17_combout;
wire fxp_functions_0_aMux_64_a0_combout;
wire fxp_functions_0_areduce_nor_18_a0_combout;
wire fxp_functions_0_areduce_nor_18_a1_combout;
wire fxp_functions_0_areduce_nor_18_a2_combout;
wire fxp_functions_0_areduce_nor_18_a3_combout;
wire fxp_functions_0_areduce_nor_18_a4_combout;
wire fxp_functions_0_areduce_nor_18_a5_combout;
wire fxp_functions_0_areduce_nor_18_a6_combout;
wire fxp_functions_0_areduce_nor_18_acombout;
wire fxp_functions_0_ai8489_a32_combout;
wire fxp_functions_0_ai8489_a33_combout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0_combout;
wire fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0_combout;
wire fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15_combout;
wire fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16_combout;
wire fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell_combout;
wire fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell_combout;
wire fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell_combout;

wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [63:0] fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus;
wire [63:0] fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus;
wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [63:0] fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [63:0] fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus;
wire [63:0] fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus;
wire [63:0] fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [63:0] fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus;
wire [143:0] fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus;
wire [19:0] fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus;

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a0_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a1_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a2_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a3_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a4_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a5_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a6_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a7_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a8_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a9_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a10_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a11_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a12_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a13_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a14_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a15_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a16_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a17_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a18_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a19_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a20_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a21_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a22_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a23_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a24_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a25_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a26_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a27_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a28_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a29_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a30_a = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA31 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA32 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA33 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA34 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA35 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA36 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA37 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA38 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA39 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA40 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA41 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA42 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA43 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA44 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA45 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA46 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA47 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA48 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA49 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA50 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA51 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA52 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA53 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA54 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA55 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA56 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA57 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA58 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA59 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA60 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA61 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA62 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_aDATAOUTA63 = fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a0_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a1_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a2_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a3_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a4_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a5_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a6_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a7_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a8_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a9_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a10_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a11_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a12_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a13_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a14_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a15_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a16_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a17_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a18_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a19_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a20_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a21_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a22_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a23_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a24_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a25_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a26_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a27_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a28_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a29_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a30_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a31_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a32_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a33_a = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA34 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA35 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA36 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA37 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA38 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA39 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA40 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA41 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA42 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA43 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA44 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA45 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA46 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA47 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA48 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA49 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA50 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA51 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA52 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA53 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA54 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA55 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA56 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA57 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA58 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA59 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA60 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA61 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA62 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_aDATAOUTA63 = fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a0_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a1_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a2_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a3_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a4_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a5_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a6_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a7_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a8_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a9_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a10_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a11_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a12_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a13_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a14_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a15_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a16_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a17_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a18_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a19_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a20_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a21_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a22_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a23_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a24_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a25_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a26_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a27_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a28_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a29_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a30_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a31_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a32_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a33_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a34_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a35_a = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA36 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA37 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA38 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA39 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA40 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA41 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA42 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA43 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA44 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA45 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA46 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA47 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA48 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA49 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA50 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA51 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA52 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA53 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA54 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA55 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA56 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA57 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA58 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA59 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA60 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA61 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA62 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_aDATAOUTA63 = fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a24_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a25_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a26_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a27_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a28_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a29_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a30_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a31_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus[19];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a30_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a31_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a32_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a33_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a34_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a35_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a36_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36_PORTBDATAOUT_bus[0];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19 = fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[19];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a0_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a1_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a2_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a3_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a4_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a5_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a6_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a7_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a8_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a9_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a10_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a11_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a12_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a13_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a14_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a15_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a16_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a17_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a18_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a19_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a20_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a21_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a22_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a23_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a24_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a25_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a26_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a27_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a28_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a29_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a30_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a31_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a32_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a33_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a34_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a35_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a36_a = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA37 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA38 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA39 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA40 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA41 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA42 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA43 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA44 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA45 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA46 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA47 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA48 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA49 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA50 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA51 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA52 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA53 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA54 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA55 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA56 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA57 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA58 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA59 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA60 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA61 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA62 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA63 = fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a0_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a1_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a2_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a3_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a4_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a5_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a6_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a7_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a8_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a9_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a10_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a11_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a12_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a13_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a14_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a15_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a16_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a17_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a18_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a19_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a20_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a21_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a22_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a23_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a24_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a25_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a26_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a27_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a28_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a29_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a30_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a31_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a32_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a33_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a34_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a35_a = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA36 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA37 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA38 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA39 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA40 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA41 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA42 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA43 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA44 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA45 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA46 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA47 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA48 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA49 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA50 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA51 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA52 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA53 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA54 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA55 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA56 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA57 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA58 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA59 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA60 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA61 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA62 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_aDATAOUTA63 = fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a0_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a1_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a2_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a3_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a4_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a5_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a6_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a7_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a8_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a9_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a10_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a11_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a12_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a13_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a14_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a15_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a16_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a17_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a18_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a19_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a20_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a21_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a22_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a23_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a24_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a25_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a26_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a27_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a28_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a29_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a30_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a31_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a32_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a33_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a34_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a35_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a36_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a37_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a38_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a39_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a40_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a41_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a42_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a43_a = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA44 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA45 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA46 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA47 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA48 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA49 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA50 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA51 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA52 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA53 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA54 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA55 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA56 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA57 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA58 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA59 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA60 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA61 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA62 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_aDATAOUTA63 = fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a = fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus[0];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a0_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[0];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a1_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[1];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a2_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[2];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a3_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[3];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a4_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[4];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a5_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[5];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a6_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[6];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a7_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[7];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a8_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[8];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a9_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[9];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a10_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[10];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a11_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[11];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a12_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[12];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a13_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[13];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a14_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[14];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a15_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[15];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a16_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[16];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a17_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[17];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a18_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[18];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a19_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[19];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a20_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[20];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a21_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[21];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a22_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[22];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a23_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[23];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a24_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[24];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a25_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[25];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a26_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[26];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a27_a = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[27];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA28 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[28];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA29 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[29];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA30 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[30];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA31 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[31];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA32 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[32];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA33 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[33];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA34 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[34];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA35 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[35];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA36 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[36];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA37 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[37];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA38 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[38];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA39 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[39];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA40 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[40];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA41 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[41];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA42 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[42];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA43 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[43];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA44 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[44];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA45 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[45];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA46 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[46];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA47 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[47];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA48 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[48];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA49 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[49];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA50 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[50];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA51 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[51];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA52 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[52];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA53 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[53];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA54 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[54];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA55 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[55];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA56 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[56];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA57 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[57];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA58 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[58];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA59 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[59];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA60 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[60];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA61 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[61];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA62 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[62];
assign fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_aDATAOUTA63 = fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus[63];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a = fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus[0];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus[0];

assign fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a = fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus[0];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus[19];

assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[0];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT1 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[1];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT2 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[2];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT3 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[3];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT4 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[4];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT5 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[5];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT6 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[6];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT7 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[7];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT8 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[8];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT9 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[9];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT10 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[10];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT11 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[11];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT12 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[12];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT13 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[13];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT14 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[14];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT15 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[15];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT16 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[16];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT17 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[17];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT18 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[18];
assign fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_aPORTBDATAOUT19 = fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus[19];

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a151_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_17_a156_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a_aq));
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a162_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a1_sumout),
	.cout(fxp_functions_0_aadd_17_a2),
	.shareout());
defparam fxp_functions_0_aadd_17_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a1.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a6_sumout),
	.cout(fxp_functions_0_aadd_17_a7),
	.shareout());
defparam fxp_functions_0_aadd_17_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a6.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a11_sumout),
	.cout(fxp_functions_0_aadd_17_a12),
	.shareout());
defparam fxp_functions_0_aadd_17_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a11.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a16_sumout),
	.cout(fxp_functions_0_aadd_17_a17),
	.shareout());
defparam fxp_functions_0_aadd_17_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a16.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a21_sumout),
	.cout(fxp_functions_0_aadd_17_a22),
	.shareout());
defparam fxp_functions_0_aadd_17_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a21.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a26_sumout),
	.cout(fxp_functions_0_aadd_17_a27),
	.shareout());
defparam fxp_functions_0_aadd_17_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a26.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a31_sumout),
	.cout(fxp_functions_0_aadd_17_a32),
	.shareout());
defparam fxp_functions_0_aadd_17_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a31.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a36_sumout),
	.cout(fxp_functions_0_aadd_17_a37),
	.shareout());
defparam fxp_functions_0_aadd_17_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a36.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a41_sumout),
	.cout(fxp_functions_0_aadd_17_a42),
	.shareout());
defparam fxp_functions_0_aadd_17_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a41.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a46_sumout),
	.cout(fxp_functions_0_aadd_17_a47),
	.shareout());
defparam fxp_functions_0_aadd_17_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a46.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a51_sumout),
	.cout(fxp_functions_0_aadd_17_a52),
	.shareout());
defparam fxp_functions_0_aadd_17_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a51.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a56_sumout),
	.cout(fxp_functions_0_aadd_17_a57),
	.shareout());
defparam fxp_functions_0_aadd_17_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a56.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a61_sumout),
	.cout(fxp_functions_0_aadd_17_a62),
	.shareout());
defparam fxp_functions_0_aadd_17_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a61.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a66_sumout),
	.cout(fxp_functions_0_aadd_17_a67),
	.shareout());
defparam fxp_functions_0_aadd_17_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a66.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a71_sumout),
	.cout(fxp_functions_0_aadd_17_a72),
	.shareout());
defparam fxp_functions_0_aadd_17_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a71.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a76_sumout),
	.cout(fxp_functions_0_aadd_17_a77),
	.shareout());
defparam fxp_functions_0_aadd_17_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a76.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a81_sumout),
	.cout(fxp_functions_0_aadd_17_a82),
	.shareout());
defparam fxp_functions_0_aadd_17_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a81.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a86_sumout),
	.cout(fxp_functions_0_aadd_17_a87),
	.shareout());
defparam fxp_functions_0_aadd_17_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a86.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a91_sumout),
	.cout(fxp_functions_0_aadd_17_a92),
	.shareout());
defparam fxp_functions_0_aadd_17_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a91.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a96_sumout),
	.cout(fxp_functions_0_aadd_17_a97),
	.shareout());
defparam fxp_functions_0_aadd_17_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a96.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a101_sumout),
	.cout(fxp_functions_0_aadd_17_a102),
	.shareout());
defparam fxp_functions_0_aadd_17_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a101.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a106_sumout),
	.cout(fxp_functions_0_aadd_17_a107),
	.shareout());
defparam fxp_functions_0_aadd_17_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a106.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a111_sumout),
	.cout(fxp_functions_0_aadd_17_a112),
	.shareout());
defparam fxp_functions_0_aadd_17_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a111.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a116_sumout),
	.cout(fxp_functions_0_aadd_17_a117),
	.shareout());
defparam fxp_functions_0_aadd_17_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a116.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a121_sumout),
	.cout(fxp_functions_0_aadd_17_a122),
	.shareout());
defparam fxp_functions_0_aadd_17_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a121.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a126_sumout),
	.cout(fxp_functions_0_aadd_17_a127),
	.shareout());
defparam fxp_functions_0_aadd_17_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a126.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a126.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a131_sumout),
	.cout(fxp_functions_0_aadd_17_a132),
	.shareout());
defparam fxp_functions_0_aadd_17_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a131.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a131.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a136_sumout),
	.cout(fxp_functions_0_aadd_17_a137),
	.shareout());
defparam fxp_functions_0_aadd_17_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a136.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a136.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a141_sumout),
	.cout(fxp_functions_0_aadd_17_a142),
	.shareout());
defparam fxp_functions_0_aadd_17_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a141.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a141.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a146_sumout),
	.cout(fxp_functions_0_aadd_17_a147),
	.shareout());
defparam fxp_functions_0_aadd_17_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a146.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a146.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a151_sumout),
	.cout(fxp_functions_0_aadd_17_a152),
	.shareout());
defparam fxp_functions_0_aadd_17_a151.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a151.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a151.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a156(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_17_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_17_a156_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_17_a156.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a156.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_17_a156.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_17_a162(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a_aq),
	.datad(!fxp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_17_a162_cout),
	.shareout());
defparam fxp_functions_0_aadd_17_a162.extended_lut = "off";
defparam fxp_functions_0_aadd_17_a162.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_17_a162.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a79_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a74_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a69_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a64_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a59_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a54_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a49_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a44_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a39_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a34_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_176_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_175_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_174_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_173_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_172_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_171_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_170_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_169_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_168_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_167_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_166_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_165_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_164_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_163_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_162_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_arShiftCount_uid26_divider_o_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq));
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_arShiftCount_uid26_divider_o_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a151_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a156_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a161_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a157),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a1_sumout),
	.cout(fxp_functions_0_aadd_13_a2),
	.shareout());
defparam fxp_functions_0_aadd_13_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a1.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a6_sumout),
	.cout(fxp_functions_0_aadd_13_a7),
	.shareout());
defparam fxp_functions_0_aadd_13_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a6.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a11_sumout),
	.cout(fxp_functions_0_aadd_13_a12),
	.shareout());
defparam fxp_functions_0_aadd_13_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a11.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a16_sumout),
	.cout(fxp_functions_0_aadd_13_a17),
	.shareout());
defparam fxp_functions_0_aadd_13_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a16.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a21_sumout),
	.cout(fxp_functions_0_aadd_13_a22),
	.shareout());
defparam fxp_functions_0_aadd_13_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a21.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a26_sumout),
	.cout(fxp_functions_0_aadd_13_a27),
	.shareout());
defparam fxp_functions_0_aadd_13_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a26.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a31_sumout),
	.cout(fxp_functions_0_aadd_13_a32),
	.shareout());
defparam fxp_functions_0_aadd_13_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a31.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a36_sumout),
	.cout(fxp_functions_0_aadd_13_a37),
	.shareout());
defparam fxp_functions_0_aadd_13_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a36.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a41_sumout),
	.cout(fxp_functions_0_aadd_13_a42),
	.shareout());
defparam fxp_functions_0_aadd_13_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a41.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a46_sumout),
	.cout(fxp_functions_0_aadd_13_a47),
	.shareout());
defparam fxp_functions_0_aadd_13_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a46.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a51_sumout),
	.cout(fxp_functions_0_aadd_13_a52),
	.shareout());
defparam fxp_functions_0_aadd_13_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a51.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a56_sumout),
	.cout(fxp_functions_0_aadd_13_a57),
	.shareout());
defparam fxp_functions_0_aadd_13_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a56.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a61_sumout),
	.cout(fxp_functions_0_aadd_13_a62),
	.shareout());
defparam fxp_functions_0_aadd_13_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a61.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a66_sumout),
	.cout(fxp_functions_0_aadd_13_a67),
	.shareout());
defparam fxp_functions_0_aadd_13_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a66.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a71_sumout),
	.cout(fxp_functions_0_aadd_13_a72),
	.shareout());
defparam fxp_functions_0_aadd_13_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a71.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a76_sumout),
	.cout(fxp_functions_0_aadd_13_a77),
	.shareout());
defparam fxp_functions_0_aadd_13_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a76.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a76.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a167),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a81_sumout),
	.cout(fxp_functions_0_aadd_13_a82),
	.shareout());
defparam fxp_functions_0_aadd_13_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a86_sumout),
	.cout(fxp_functions_0_aadd_13_a87),
	.shareout());
defparam fxp_functions_0_aadd_13_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a86.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a91_sumout),
	.cout(fxp_functions_0_aadd_13_a92),
	.shareout());
defparam fxp_functions_0_aadd_13_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a91.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a96_sumout),
	.cout(fxp_functions_0_aadd_13_a97),
	.shareout());
defparam fxp_functions_0_aadd_13_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a96.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a101_sumout),
	.cout(fxp_functions_0_aadd_13_a102),
	.shareout());
defparam fxp_functions_0_aadd_13_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a101.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a106_sumout),
	.cout(fxp_functions_0_aadd_13_a107),
	.shareout());
defparam fxp_functions_0_aadd_13_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a106.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a111_sumout),
	.cout(fxp_functions_0_aadd_13_a112),
	.shareout());
defparam fxp_functions_0_aadd_13_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a111.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a116_sumout),
	.cout(fxp_functions_0_aadd_13_a117),
	.shareout());
defparam fxp_functions_0_aadd_13_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a116.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a121_sumout),
	.cout(fxp_functions_0_aadd_13_a122),
	.shareout());
defparam fxp_functions_0_aadd_13_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a121.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a126_sumout),
	.cout(fxp_functions_0_aadd_13_a127),
	.shareout());
defparam fxp_functions_0_aadd_13_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a126.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a126.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a131_sumout),
	.cout(fxp_functions_0_aadd_13_a132),
	.shareout());
defparam fxp_functions_0_aadd_13_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a131.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a131.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a136_sumout),
	.cout(fxp_functions_0_aadd_13_a137),
	.shareout());
defparam fxp_functions_0_aadd_13_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a136.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a136.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a141_sumout),
	.cout(fxp_functions_0_aadd_13_a142),
	.shareout());
defparam fxp_functions_0_aadd_13_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a141.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a141.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a146_sumout),
	.cout(fxp_functions_0_aadd_13_a147),
	.shareout());
defparam fxp_functions_0_aadd_13_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a146.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a146.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a151_sumout),
	.cout(fxp_functions_0_aadd_13_a152),
	.shareout());
defparam fxp_functions_0_aadd_13_a151.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a151.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a151.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a156(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a156_sumout),
	.cout(fxp_functions_0_aadd_13_a157),
	.shareout());
defparam fxp_functions_0_aadd_13_a156.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a156.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a156.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_13_a166_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a161(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a161_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_13_a161.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a161.lut_mask = 64'h0000000000000F0F;
defparam fxp_functions_0_aadd_13_a161.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a166(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a172_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_13_a166_sumout),
	.cout(fxp_functions_0_aadd_13_a167),
	.shareout());
defparam fxp_functions_0_aadd_13_a166.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a166.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a166.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai8103_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mac fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.ax_width = 15;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.ay_scan_in_width = 16;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.result_a_width = 31;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.signed_may = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_DSP0.use_chainadder = "false";

fourteennm_mac fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx({fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a_aq}),
	.by({gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a_aq}),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.ay_scan_in_width = 15;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.bx_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.bx_width = 18;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.by_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.by_width = 15;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.operation_mode = "m18x18_sumof2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.result_a_width = 34;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.signed_max = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_DSP0.use_chainadder = "false";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 5;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 28;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 29;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist11_r_uid72_zcount_uid9_divider_q_32_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 6;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mac fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a_aq,
fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a_aq,fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.ay_scan_in_width = 18;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.result_a_width = 36;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.signed_max = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_DSP0.use_chainadder = "false";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a172(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a177_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a172_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a172.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a172.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a172.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_21_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a177(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a182_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a177_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a177.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a177.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a177.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_15_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai8126_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai8126_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai8126_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a20_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a22_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a23_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a24_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a25_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a26_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a27_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a28_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a29_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a30_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a31_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_ai6816_a32_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a_aq));
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_10_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_9_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq));
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a182(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a187_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a182_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a182.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a182.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a182.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_17_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a_aq));
defparam fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a_aq));
defparam fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a162),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a1_sumout),
	.cout(fxp_functions_0_aadd_12_a2),
	.shareout());
defparam fxp_functions_0_aadd_12_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a1.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a6_sumout),
	.cout(fxp_functions_0_aadd_12_a7),
	.shareout());
defparam fxp_functions_0_aadd_12_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a6.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a11_sumout),
	.cout(fxp_functions_0_aadd_12_a12),
	.shareout());
defparam fxp_functions_0_aadd_12_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a11.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a16_sumout),
	.cout(fxp_functions_0_aadd_12_a17),
	.shareout());
defparam fxp_functions_0_aadd_12_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a21_sumout),
	.cout(fxp_functions_0_aadd_12_a22),
	.shareout());
defparam fxp_functions_0_aadd_12_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a21.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a26_sumout),
	.cout(fxp_functions_0_aadd_12_a27),
	.shareout());
defparam fxp_functions_0_aadd_12_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a26.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a31_sumout),
	.cout(fxp_functions_0_aadd_12_a32),
	.shareout());
defparam fxp_functions_0_aadd_12_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a31.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a29_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a36_sumout),
	.cout(fxp_functions_0_aadd_12_a37),
	.shareout());
defparam fxp_functions_0_aadd_12_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a36.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a41(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a30_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a41_sumout),
	.cout(fxp_functions_0_aadd_12_a42),
	.shareout());
defparam fxp_functions_0_aadd_12_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a41.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a46(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a31_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a46_sumout),
	.cout(fxp_functions_0_aadd_12_a47),
	.shareout());
defparam fxp_functions_0_aadd_12_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a46.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a51(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a32_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a51_sumout),
	.cout(fxp_functions_0_aadd_12_a52),
	.shareout());
defparam fxp_functions_0_aadd_12_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a51.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a56(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a33_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a56_sumout),
	.cout(fxp_functions_0_aadd_12_a57),
	.shareout());
defparam fxp_functions_0_aadd_12_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a56.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a61(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a34_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a61_sumout),
	.cout(fxp_functions_0_aadd_12_a62),
	.shareout());
defparam fxp_functions_0_aadd_12_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a61.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a66(
	.dataa(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a35_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a66_sumout),
	.cout(fxp_functions_0_aadd_12_a67),
	.shareout());
defparam fxp_functions_0_aadd_12_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a66.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_12_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a36_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a71_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_12_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a71.lut_mask = 64'h0000000000000FF0;
defparam fxp_functions_0_aadd_12_a71.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a167_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a76_sumout),
	.cout(fxp_functions_0_aadd_12_a77),
	.shareout());
defparam fxp_functions_0_aadd_12_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a76.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a81_sumout),
	.cout(fxp_functions_0_aadd_12_a82),
	.shareout());
defparam fxp_functions_0_aadd_12_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a86_sumout),
	.cout(fxp_functions_0_aadd_12_a87),
	.shareout());
defparam fxp_functions_0_aadd_12_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a86.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a91_sumout),
	.cout(fxp_functions_0_aadd_12_a92),
	.shareout());
defparam fxp_functions_0_aadd_12_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a91.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a96_sumout),
	.cout(fxp_functions_0_aadd_12_a97),
	.shareout());
defparam fxp_functions_0_aadd_12_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a96.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a101_sumout),
	.cout(fxp_functions_0_aadd_12_a102),
	.shareout());
defparam fxp_functions_0_aadd_12_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a101.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a106_sumout),
	.cout(fxp_functions_0_aadd_12_a107),
	.shareout());
defparam fxp_functions_0_aadd_12_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a106.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a111_sumout),
	.cout(fxp_functions_0_aadd_12_a112),
	.shareout());
defparam fxp_functions_0_aadd_12_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a111.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a116_sumout),
	.cout(fxp_functions_0_aadd_12_a117),
	.shareout());
defparam fxp_functions_0_aadd_12_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a116.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a121_sumout),
	.cout(fxp_functions_0_aadd_12_a122),
	.shareout());
defparam fxp_functions_0_aadd_12_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a121.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a126_sumout),
	.cout(fxp_functions_0_aadd_12_a127),
	.shareout());
defparam fxp_functions_0_aadd_12_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a126.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a126.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a131_sumout),
	.cout(fxp_functions_0_aadd_12_a132),
	.shareout());
defparam fxp_functions_0_aadd_12_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a131.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a131.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a136_sumout),
	.cout(fxp_functions_0_aadd_12_a137),
	.shareout());
defparam fxp_functions_0_aadd_12_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a136.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a136.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a141_sumout),
	.cout(fxp_functions_0_aadd_12_a142),
	.shareout());
defparam fxp_functions_0_aadd_12_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a141.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a141.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a146_sumout),
	.cout(fxp_functions_0_aadd_12_a147),
	.shareout());
defparam fxp_functions_0_aadd_12_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a146.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a146.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a151_sumout),
	.cout(fxp_functions_0_aadd_12_a152),
	.shareout());
defparam fxp_functions_0_aadd_12_a151.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a151.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a151.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a156(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a156_sumout),
	.cout(fxp_functions_0_aadd_12_a157),
	.shareout());
defparam fxp_functions_0_aadd_12_a156.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a156.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a156.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a161(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a157),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_12_a161_sumout),
	.cout(fxp_functions_0_aadd_12_a162),
	.shareout());
defparam fxp_functions_0_aadd_12_a161.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a161.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a161.shared_arith = "off";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai3244_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a_aq));
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_8_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a_aq));
defparam fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist12_vCount_uid53_zCount_uid9_divider_q_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a187(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a192_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a187_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a187.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a187.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a187.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_7_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a_aq));
defparam fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist13_vCount_uid47_zCount_uid9_divider_q_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a(
	.clk(clk),
	.d(fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a_aq));
defparam fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist14_vCount_uid41_zCount_uid9_divider_q_3_delay_0_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_bit_number = 18;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama18";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai1590_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_bit_number = 19;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama19";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_bit_number = 20;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama20";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_bit_number = 21;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama21";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_bit_number = 22;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama22";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.first_bit_number = 23;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama23";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama23.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.first_bit_number = 24;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama24";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama24.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.first_bit_number = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama25";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama25.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.first_bit_number = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama26";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama26.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.first_bit_number = 27;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama27";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama27.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.first_bit_number = 28;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama28";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama28.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.first_bit_number = 29;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama29";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama29.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.first_bit_number = 30;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama30";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama30.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.first_bit_number = 31;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama31";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama31.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_bit_number = 22;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_bit_number = 22;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mem_init0 = "066AB61E32A90E12AC3194C06A9F1588D31D60D3CA05797D7D3319AF45E68B90";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_bit_number = 23;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_bit_number = 23;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mem_init0 = "01E66D4B5B31F1F19A9AD8FFE64A59F7C9567FC96C032D8329CEAE65834653B8";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_bit_number = 24;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_bit_number = 24;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mem_init0 = "001E1CC6C96B555AD3231F001E3934AA92678038DAAA4E00E4AB301CAA79C920";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_bit_number = 25;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_bit_number = 25;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mem_init0 = "0001FC3E38E7333649694AAAAB5259331C780007C666DAAAB6CC3FFC66D56DC0";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a28_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_bit_number = 26;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_bit_number = 26;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mem_init0 = "AAAAA954AD4A5A5B6DB26CCCCC639E3C1F8000003E1E3999925A9556B4998E00";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a29_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_bit_number = 27;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_bit_number = 27;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mem_init0 = "666664CD9B26C936DB6925A5A5294A954AAAAAAAAB54AD2D2493266738E1F000";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a30_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_bit_number = 28;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_bit_number = 28;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mem_init0 = "1E1E1C3C78E1C70E38E71C639CE7398CC666666666CD9B6492496D2D6A54AAAA";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a31_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_first_bit_number = 29;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_first_bit_number = 29;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a29.mem_init0 = "01FE03FC07E03F01F81F03E07C1F0783C1E1E1E1E1C3871C71C71CE319CC6666";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_first_bit_number = 30;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_first_bit_number = 30;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a30.mem_init0 = "0001FFFC001FFF0007FF001FFC00FF803FE01FE01FC07F03F03F03E0F83C1E1E";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_first_bit_number = 31;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_first_bit_number = 31;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a31.mem_init0 = "00000003FFFFFF000000FFFFFC00007FFFE0001FFFC000FFF000FFE007FC01FE";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_first_bit_number = 32;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_first_bit_number = 32;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a32.mem_init0 = "00000000000000FFFFFFFFFFFC000000001FFFFFFFC000000FFFFFE00003FFFE";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_first_bit_number = 33;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_first_bit_number = 33;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a33.mem_init0 = "00000000000000000000000003FFFFFFFFFFFFFFFFC000000000001FFFFFFFFE";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_first_bit_number = 34;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_first_bit_number = 34;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a34.mem_init0 = "0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFE";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_first_bit_number = 35;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_first_bit_number = 35;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a35.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_first_bit_number = 36;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_first_bit_number = 36;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a36.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000001";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_bit_number = 16;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama16";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq}),
	.portaaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.address_width = 5;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.data_width = 1;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_address = 0;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_bit_number = 17;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.init_file = "none";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.last_address = 25;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_depth = 26;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_name = "fxp_functions_0|redist21_in_rsrvd_fix_numerator_29_mem_dmem|auto_generated|altera_syncram_impl1|lutrama17";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_width = 32;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "0470BC98F923B85E09A97FCDBCB76F9C28B802296EB55F2960B1F60944A9B0A2";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a167(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a172_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_12_a167_cout),
	.shareout());
defparam fxp_functions_0_aadd_12_a167.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a167.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a167.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "217791106142C56123A4AE6810DE329762D0C56704A19A58E3D4FD054DD09A40";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "0A5A2378A01E930CFF91A2F37C6D4A9E91C21BA83D0EC37B464FBDF40058B930";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "1642C135F9FB9D1203594DF9A6556D612D85844E39C8156B36AA8EDED520F410";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "A254BB9A45088C8B86A295D90C8DC79A87847BE48A0633A8EBCE2A30A4331C5C";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "2EC827A24F00BB42A0710A8455D72F4B4224B1BF4040B53272CB15A16F5F20F0";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "088F555AAD623744BB71BF8694002A14C54B4A5C0C55977FCD0F26699D0BDA78";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "6F58C8AF91B22787FE8125FBB7220A49D8673D3522D5E2B53D27950BA95B8F50";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "2E62EC5A4201BF0CF9438B4654FAF3B2DD7E68CD4844E234845B9EA80234BF2A";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "08D00DB84181E904E2143DE88A1D48BF0E9D445FC9C66274C43268A2885CCB82";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "1EF8A64A6A4C303310E70B68F20C7F328AC28402D262ED1596411862368C776A";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "04DBFB1B26870C7AA13472616CADE29FCCD8AA4103E4D5CB64D891FD64089746";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "0266EE222D6474566A1A30A90A663AB8B0CEA8C08F0D8AEA3631CA75D8656686";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "AB7E4EB80DC09F5780C72DC659E2B89BE6A2EDC051C5C8A6B139469FBFC506CE";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "00B2E80A7FB1C42088BACBF5381E6C8C4345F70CF91818CB321AA7C42A81601E";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "444A6117C71D8A36BEB06B3561987C49B24E244B43141259640C438A5565F0BE";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "282DCF5E8209AEB36E34361B90F16D2A4AAC55FE0E80D05E8B364DC8EEF250D4";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_bit_number = 21;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_bit_number = 21;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mem_init0 = "1AB0259E5404CE641B32BEA0A05F334978E7DB7BD1086BE444B6AD81393603D4";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a22_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai3159_a23_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a_aq));
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a192(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a197_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a192_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a192.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a192.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a192.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_6_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a(
	.clk(clk),
	.d(denominator[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a(
	.clk(clk),
	.d(denominator[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a(
	.clk(clk),
	.d(denominator[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a(
	.clk(clk),
	.d(denominator[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a(
	.clk(clk),
	.d(denominator[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a(
	.clk(clk),
	.d(denominator[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a(
	.clk(clk),
	.d(denominator[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a(
	.clk(clk),
	.d(denominator[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a(
	.clk(clk),
	.d(denominator[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a(
	.clk(clk),
	.d(denominator[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a(
	.clk(clk),
	.d(denominator[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a(
	.clk(clk),
	.d(denominator[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a(
	.clk(clk),
	.d(denominator[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a(
	.clk(clk),
	.d(denominator[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a(
	.clk(clk),
	.d(denominator[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a(
	.clk(clk),
	.d(denominator[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_19_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a2_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a1(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a1_sumout),
	.cout(fxp_functions_0_aadd_9_a2),
	.shareout());
defparam fxp_functions_0_aadd_9_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a1.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a6(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a6_sumout),
	.cout(fxp_functions_0_aadd_9_a7),
	.shareout());
defparam fxp_functions_0_aadd_9_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a6.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a11(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a11_sumout),
	.cout(fxp_functions_0_aadd_9_a12),
	.shareout());
defparam fxp_functions_0_aadd_9_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a11.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a16(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a16_sumout),
	.cout(fxp_functions_0_aadd_9_a17),
	.shareout());
defparam fxp_functions_0_aadd_9_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a16.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a21(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a21_sumout),
	.cout(fxp_functions_0_aadd_9_a22),
	.shareout());
defparam fxp_functions_0_aadd_9_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a21.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a26(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a26_sumout),
	.cout(fxp_functions_0_aadd_9_a27),
	.shareout());
defparam fxp_functions_0_aadd_9_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a26.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a31(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a31_sumout),
	.cout(fxp_functions_0_aadd_9_a32),
	.shareout());
defparam fxp_functions_0_aadd_9_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a31.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a36_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_9_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a36.lut_mask = 64'h0000000000000FF0;
defparam fxp_functions_0_aadd_9_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a41_sumout),
	.cout(fxp_functions_0_aadd_9_a42),
	.shareout());
defparam fxp_functions_0_aadd_9_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a41.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a41.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "60B4BAC9BD0C8861A48C7921276D712D43EB4C304A045656B0FA50CB04801040";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a172(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a177_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_12_a172_cout),
	.shareout());
defparam fxp_functions_0_aadd_12_a172.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a172.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a172.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a46_sumout),
	.cout(fxp_functions_0_aadd_9_a47),
	.shareout());
defparam fxp_functions_0_aadd_9_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a46.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a51_sumout),
	.cout(fxp_functions_0_aadd_9_a52),
	.shareout());
defparam fxp_functions_0_aadd_9_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a51.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a56_sumout),
	.cout(fxp_functions_0_aadd_9_a57),
	.shareout());
defparam fxp_functions_0_aadd_9_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a56.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a61_sumout),
	.cout(fxp_functions_0_aadd_9_a62),
	.shareout());
defparam fxp_functions_0_aadd_9_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a61.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a66_sumout),
	.cout(fxp_functions_0_aadd_9_a67),
	.shareout());
defparam fxp_functions_0_aadd_9_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a66.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a71_sumout),
	.cout(fxp_functions_0_aadd_9_a72),
	.shareout());
defparam fxp_functions_0_aadd_9_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a71.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a76_sumout),
	.cout(fxp_functions_0_aadd_9_a77),
	.shareout());
defparam fxp_functions_0_aadd_9_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a76.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a81_sumout),
	.cout(fxp_functions_0_aadd_9_a82),
	.shareout());
defparam fxp_functions_0_aadd_9_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a86(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a86_sumout),
	.cout(fxp_functions_0_aadd_9_a87),
	.shareout());
defparam fxp_functions_0_aadd_9_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a86.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a91(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a91_sumout),
	.cout(fxp_functions_0_aadd_9_a92),
	.shareout());
defparam fxp_functions_0_aadd_9_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a91.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a96(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a96_sumout),
	.cout(fxp_functions_0_aadd_9_a97),
	.shareout());
defparam fxp_functions_0_aadd_9_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a96.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a101(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a101_sumout),
	.cout(fxp_functions_0_aadd_9_a102),
	.shareout());
defparam fxp_functions_0_aadd_9_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a101.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a106(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a106_sumout),
	.cout(fxp_functions_0_aadd_9_a107),
	.shareout());
defparam fxp_functions_0_aadd_9_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a106.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a111(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a111_sumout),
	.cout(fxp_functions_0_aadd_9_a112),
	.shareout());
defparam fxp_functions_0_aadd_9_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a111.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a116(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a116_sumout),
	.cout(fxp_functions_0_aadd_9_a117),
	.shareout());
defparam fxp_functions_0_aadd_9_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a116.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a121(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a121_sumout),
	.cout(fxp_functions_0_aadd_9_a122),
	.shareout());
defparam fxp_functions_0_aadd_9_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a121.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a126(
	.dataa(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a126_sumout),
	.cout(fxp_functions_0_aadd_9_a127),
	.shareout());
defparam fxp_functions_0_aadd_9_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a126.lut_mask = 64'h0000000005055A5A;
defparam fxp_functions_0_aadd_9_a126.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a(
	.clk(clk),
	.d(denominator[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a(
	.clk(clk),
	.d(denominator[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a(
	.clk(clk),
	.d(denominator[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a(
	.clk(clk),
	.d(denominator[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a(
	.clk(clk),
	.d(denominator[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a(
	.clk(clk),
	.d(denominator[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a(
	.clk(clk),
	.d(denominator[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a(
	.clk(clk),
	.d(denominator[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a(
	.clk(clk),
	.d(denominator[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a(
	.clk(clk),
	.d(denominator[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a(
	.clk(clk),
	.d(denominator[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a(
	.clk(clk),
	.d(denominator[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a(
	.clk(clk),
	.d(denominator[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a(
	.clk(clk),
	.d(denominator[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a(
	.clk(clk),
	.d(denominator[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a197(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a202_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a197_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a197.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a197.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a197.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_0_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_0_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_0_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_0_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a(
	.clk(clk),
	.d(numerator[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a(
	.clk(clk),
	.d(numerator[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a(
	.clk(clk),
	.d(numerator[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a(
	.clk(clk),
	.d(numerator[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a(
	.clk(clk),
	.d(numerator[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a(
	.clk(clk),
	.d(numerator[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a(
	.clk(clk),
	.d(numerator[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a(
	.clk(clk),
	.d(numerator[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a(
	.clk(clk),
	.d(numerator[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a(
	.clk(clk),
	.d(numerator[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a(
	.clk(clk),
	.d(numerator[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a(
	.clk(clk),
	.d(numerator[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a(
	.clk(clk),
	.d(numerator[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a(
	.clk(clk),
	.d(numerator[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a3_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a(
	.clk(clk),
	.d(numerator[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a(
	.clk(clk),
	.d(numerator[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a(
	.clk(clk),
	.d(numerator[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a(
	.clk(clk),
	.d(numerator[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a(
	.clk(clk),
	.d(numerator[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a(
	.clk(clk),
	.d(numerator[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a(
	.clk(clk),
	.d(numerator[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a(
	.clk(clk),
	.d(numerator[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a(
	.clk(clk),
	.d(numerator[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a(
	.clk(clk),
	.d(numerator[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a(
	.clk(clk),
	.d(numerator[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a(
	.clk(clk),
	.d(numerator[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a(
	.clk(clk),
	.d(numerator[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a(
	.clk(clk),
	.d(numerator[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a(
	.clk(clk),
	.d(numerator[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a(
	.clk(clk),
	.d(numerator[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a(
	.clk(clk),
	.d(numerator[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a(
	.clk(clk),
	.d(numerator[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a131_sumout),
	.cout(fxp_functions_0_aadd_9_a132),
	.shareout());
defparam fxp_functions_0_aadd_9_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a131.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a131.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "F7B1E4FB195AD798F9D1C2999D54FC755D4C77E6CC6DAED8DB670175398A56BB";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a177(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_12_a182_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_12_a177_cout),
	.shareout());
defparam fxp_functions_0_aadd_12_a177.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a177.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a177.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a202(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a207_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a202_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a202.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a202.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a202.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_2_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a4_a_a0_a.power_up = "dont_care";

fourteennm_mac fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx({fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.by({gnd,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq,
fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq,fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.ay_scan_in_width = 18;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.bx_clock = "0";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.bx_width = 18;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.by_clock = "0";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.by_width = 18;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.operation_mode = "m18x18_sumof2";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.result_a_width = 37;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.signed_mbx = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_mac fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq,
fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq,fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.ax_width = 18;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.ay_scan_in_width = 18;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.result_a_width = 36;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.signed_may = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai6102_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fxp_functions_0|redist2_yaddr_uid19_divider_merged_bit_select_b_22_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a136_sumout),
	.cout(fxp_functions_0_aadd_9_a137),
	.shareout());
defparam fxp_functions_0_aadd_9_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a136.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a136.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "00808F9C7BA46800218E9148DBE52F878981865D4B00513EE206486EDEA18304";

fourteennm_lcell_comb fxp_functions_0_aadd_12_a182(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a_aq),
	.datad(!fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_12_a182_cout),
	.shareout());
defparam fxp_functions_0_aadd_12_a182.extended_lut = "off";
defparam fxp_functions_0_aadd_12_a182.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_12_a182.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a207(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a212_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a207_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a207.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a207.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a207.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a5_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_13_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a141_sumout),
	.cout(fxp_functions_0_aadd_9_a142),
	.shareout());
defparam fxp_functions_0_aadd_9_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a141.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a141.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_9_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist7_os_uid148_pT3_uid103_invPolyEval_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a7_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a5_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a3_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a1_a_aq,fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC0_uid74_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fxp_functions_0|memoryC0_uid74_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 38;
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC0_uid74_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "33B9CCB77751D995B87B287B2AD7FDF1142E71A7AACD2A930F158D3B65B34ED8";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a212(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a217_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a212_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a212.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a212.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a212.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a6_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a136_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a141_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_8_a146_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a_aq));
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai6114_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai6114_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai6114_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a152_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_9_a146_sumout),
	.cout(fxp_functions_0_aadd_9_a147),
	.shareout());
defparam fxp_functions_0_aadd_9_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a146.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a146.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a217(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a222_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a217_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a217.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a217.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a217.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a7_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a1_sumout),
	.cout(fxp_functions_0_aadd_8_a2),
	.shareout());
defparam fxp_functions_0_aadd_8_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a1.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a6_sumout),
	.cout(fxp_functions_0_aadd_8_a7),
	.shareout());
defparam fxp_functions_0_aadd_8_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a6.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a11_sumout),
	.cout(fxp_functions_0_aadd_8_a12),
	.shareout());
defparam fxp_functions_0_aadd_8_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a11.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a16_sumout),
	.cout(fxp_functions_0_aadd_8_a17),
	.shareout());
defparam fxp_functions_0_aadd_8_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a21_sumout),
	.cout(fxp_functions_0_aadd_8_a22),
	.shareout());
defparam fxp_functions_0_aadd_8_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a21.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a26_sumout),
	.cout(fxp_functions_0_aadd_8_a27),
	.shareout());
defparam fxp_functions_0_aadd_8_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a26.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a31_sumout),
	.cout(fxp_functions_0_aadd_8_a32),
	.shareout());
defparam fxp_functions_0_aadd_8_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a31.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a36_sumout),
	.cout(fxp_functions_0_aadd_8_a37),
	.shareout());
defparam fxp_functions_0_aadd_8_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a36.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a41_sumout),
	.cout(fxp_functions_0_aadd_8_a42),
	.shareout());
defparam fxp_functions_0_aadd_8_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a41.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a46_sumout),
	.cout(fxp_functions_0_aadd_8_a47),
	.shareout());
defparam fxp_functions_0_aadd_8_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a46.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a51_sumout),
	.cout(fxp_functions_0_aadd_8_a52),
	.shareout());
defparam fxp_functions_0_aadd_8_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a51.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a56_sumout),
	.cout(fxp_functions_0_aadd_8_a57),
	.shareout());
defparam fxp_functions_0_aadd_8_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a56.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a61_sumout),
	.cout(fxp_functions_0_aadd_8_a62),
	.shareout());
defparam fxp_functions_0_aadd_8_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a61.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a66_sumout),
	.cout(fxp_functions_0_aadd_8_a67),
	.shareout());
defparam fxp_functions_0_aadd_8_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a66.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a71_sumout),
	.cout(fxp_functions_0_aadd_8_a72),
	.shareout());
defparam fxp_functions_0_aadd_8_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a71.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a76_sumout),
	.cout(fxp_functions_0_aadd_8_a77),
	.shareout());
defparam fxp_functions_0_aadd_8_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a76.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a81_sumout),
	.cout(fxp_functions_0_aadd_8_a82),
	.shareout());
defparam fxp_functions_0_aadd_8_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a81.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a86_sumout),
	.cout(fxp_functions_0_aadd_8_a87),
	.shareout());
defparam fxp_functions_0_aadd_8_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a86.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a91_sumout),
	.cout(fxp_functions_0_aadd_8_a92),
	.shareout());
defparam fxp_functions_0_aadd_8_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a91.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a96_sumout),
	.cout(fxp_functions_0_aadd_8_a97),
	.shareout());
defparam fxp_functions_0_aadd_8_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a96.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a101_sumout),
	.cout(fxp_functions_0_aadd_8_a102),
	.shareout());
defparam fxp_functions_0_aadd_8_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a101.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a21_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a106_sumout),
	.cout(fxp_functions_0_aadd_8_a107),
	.shareout());
defparam fxp_functions_0_aadd_8_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a106.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_8_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a111(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a22_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a111_sumout),
	.cout(fxp_functions_0_aadd_8_a112),
	.shareout());
defparam fxp_functions_0_aadd_8_a111.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a111.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a111.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a116(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a23_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a116_sumout),
	.cout(fxp_functions_0_aadd_8_a117),
	.shareout());
defparam fxp_functions_0_aadd_8_a116.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a116.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a116.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a121(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a24_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a121_sumout),
	.cout(fxp_functions_0_aadd_8_a122),
	.shareout());
defparam fxp_functions_0_aadd_8_a121.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a121.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a121.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a126(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a25_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a126_sumout),
	.cout(fxp_functions_0_aadd_8_a127),
	.shareout());
defparam fxp_functions_0_aadd_8_a126.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a126.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a126.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a131(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a26_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a131_sumout),
	.cout(fxp_functions_0_aadd_8_a132),
	.shareout());
defparam fxp_functions_0_aadd_8_a131.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a131.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a131.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a136(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a27_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a136_sumout),
	.cout(fxp_functions_0_aadd_8_a137),
	.shareout());
defparam fxp_functions_0_aadd_8_a136.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a136.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_8_a136.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a141(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a141_sumout),
	.cout(fxp_functions_0_aadd_8_a142),
	.shareout());
defparam fxp_functions_0_aadd_8_a141.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a141.lut_mask = 64'h0000000011116666;
defparam fxp_functions_0_aadd_8_a141.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_8_a146(
	.dataa(!fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq),
	.datab(!fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a28_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_8_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_8_a146_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_8_a146.extended_lut = "off";
defparam fxp_functions_0_aadd_8_a146.lut_mask = 64'h0000000000006666;
defparam fxp_functions_0_aadd_8_a146.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_14_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a152(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a157_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a152_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a152.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a152.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a152.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a222(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a227_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a222_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a222.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a222.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a222.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a8_a_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai1992_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_bit_number = 16;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama16";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_bit_number = 17;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama17";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_bit_number = 18;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama18";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_bit_number = 19;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama19";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_bit_number = 20;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama20";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_bit_number = 21;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama21";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_bit_number = 22;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama22";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.mixed_port_feed_through_mode = "dont care";

fourteennm_mac fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a_aq,
fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a_aq,fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.ax_width = 23;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.ay_scan_in_width = 21;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.operation_mode = "m27x27";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.result_a_width = 44;
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "06CADCAA26E1D8F1A33773BFBBBBFF7A545C267168534FA423A66DEE2F1F1920";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "96FCABD508F2FE555FFA8B1395A0D4B3368691B10544A01AC12DC431E0DB5E6E";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "169771557E1699BA59194BAD7F0D213FF9DA9B053A10E9F5C72A5042861E3035";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "31C43729E43144D8D614F515822625C800A0073E10960D170083013A40C5944C";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "5071C41DE0ABE725028CC48DCEDEA085BC5FA554E6B950C7C397816007FF07D4";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "51C3807CCDCDEFA0C21E57C6596ECBD1A8EAC6065F02E5F44EAB8EC28CB821DC";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "776CFB7F20F752AB3A2179B6264953C09248BC052873AAA5FB073DF484D62CC6";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "6147A818B49D928D322738D40C6AF738483D7618CA1B204C0E0404F5E64F0ABC";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "D1CE01DAC66F809B2EFDA9D00B49E9FCD26ECD8B2546F6BDED6FA287FAB70914";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "57F91099ADF4384BFA4366A194F7F6CD3656D69E1EA1DCDB5707FFFFC264CFB8";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "B885F51863F97DE521197948F7D550B53D5CCD9733BFEE8F3BC28C5183932678";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "93653F818667CD92AE253A2FA7CCCF2D842EA5FCB46AA063CE2B21A8FC961F30";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "CD0D843C25A44A921725DF29F4F0F3044A39EB0867E660A2E27F0710559F334A";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "EB088681669932662F98E86C29EE12D848DC839CDE7879506FC4BDF566CF87E0";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "F25B872B18D4FCAE357EA7BBCBF5E6146741883E10F70912571B5AC01E8CE36E";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "FC6D2D6700E6AA61C6559FCD5806AE19206B8D7F4F5059B33AE842111061D802";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "FF8E364A55AD99E007992AA4C7F8CB4B1F8D24FF95306C8C560D3CB1B0A142F6";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "FFF038739936D2B552B4999C3FFF0C6DAAA49C0019A5247F9B5B00DB70CB3CAE";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "55556AD6B4924993318C787C00000F8E3336D6AAB4931C001C6DAA48F0F2559E";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "9999B364D92492DA5AD6AD56AAAAA55A96924D998C70FC001F8E336D5A56CC7E";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "E1E1C3871E38E31C6318CE673333366CDB2496D2D6A556AAB55A96DB3631C3FE";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_first_bit_number = 21;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_first_bit_number = 21;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a21.mem_init0 = "FE01FC07E03F03E07C1F0F87C3C3C78F1C38E71CE73998CCD99324925B5A9554";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_first_bit_number = 22;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_first_bit_number = 22;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a22.mem_init0 = "FFFE0007FFC003FF801FF007FC03F80FE03F07E0F83E1F0F1E1C38E39C631998";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_first_bit_number = 23;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_first_bit_number = 23;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a23.mem_init0 = "FFFFFFF8000003FFFFE00007FFFC000FFFC007FF003FE00FE01FC0FC1F83E1E0";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_first_bit_number = 24;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_first_bit_number = 24;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a24.mem_init0 = "FFFFFFFFFFFFFC0000000007FFFFFFF0000007FFFFC0000FFFE000FFE003FE00";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_first_bit_number = 25;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_first_bit_number = 25;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a25.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFF800000000000007FFFFFFFFF0000000FFFFFC0000";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_first_bit_number = 26;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_first_bit_number = 26;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a26.mem_init0 = "00000000000000000000000000000000000007FFFFFFFFFFFFFFFF0000000000";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_first_bit_number = 27;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_first_bit_number = 27;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a27.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000";

fourteennm_ram_block fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a7_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a5_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a3_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a1_a_aq,fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC1_uid77_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.logical_ram_name = "fxp_functions_0|memoryC1_uid77_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_first_bit_number = 28;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_a_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_first_bit_number = 28;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.port_b_logical_ram_width = 29;
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC1_uid77_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a28.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 2;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 3;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 4;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist5_yaddr_uid19_divider_merged_bit_select_c_17_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 23;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_q_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a157(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a162_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a157_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a157.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a157.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a157.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a227(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_13_a232_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a227_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a227.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a227.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a227.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a9_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_20_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_3_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a162(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a167_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a162_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a162.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a162.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a162.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_13_a232(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_13_a232_cout),
	.shareout());
defparam fxp_functions_0_aadd_13_a232.extended_lut = "off";
defparam fxp_functions_0_aadd_13_a232.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_13_a232.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a10_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai1997_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_2_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aadd_7_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a_aq));
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_2_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a167(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_9_a172_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a167_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a167.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a167.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a167.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a11_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a1_sumout),
	.cout(fxp_functions_0_aadd_7_a2),
	.shareout());
defparam fxp_functions_0_aadd_7_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a1.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a6_sumout),
	.cout(fxp_functions_0_aadd_7_a7),
	.shareout());
defparam fxp_functions_0_aadd_7_a6.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a6.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a11_sumout),
	.cout(fxp_functions_0_aadd_7_a12),
	.shareout());
defparam fxp_functions_0_aadd_7_a11.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a11.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a16_sumout),
	.cout(fxp_functions_0_aadd_7_a17),
	.shareout());
defparam fxp_functions_0_aadd_7_a16.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a16.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a21_sumout),
	.cout(fxp_functions_0_aadd_7_a22),
	.shareout());
defparam fxp_functions_0_aadd_7_a21.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a21.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a26_sumout),
	.cout(fxp_functions_0_aadd_7_a27),
	.shareout());
defparam fxp_functions_0_aadd_7_a26.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a26.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a31_sumout),
	.cout(fxp_functions_0_aadd_7_a32),
	.shareout());
defparam fxp_functions_0_aadd_7_a31.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a31.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a36_sumout),
	.cout(fxp_functions_0_aadd_7_a37),
	.shareout());
defparam fxp_functions_0_aadd_7_a36.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a36.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a41_sumout),
	.cout(fxp_functions_0_aadd_7_a42),
	.shareout());
defparam fxp_functions_0_aadd_7_a41.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a41.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a46_sumout),
	.cout(fxp_functions_0_aadd_7_a47),
	.shareout());
defparam fxp_functions_0_aadd_7_a46.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a46.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a51_sumout),
	.cout(fxp_functions_0_aadd_7_a52),
	.shareout());
defparam fxp_functions_0_aadd_7_a51.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a51.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a56_sumout),
	.cout(fxp_functions_0_aadd_7_a57),
	.shareout());
defparam fxp_functions_0_aadd_7_a56.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a56.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_7_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a61(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a61_sumout),
	.cout(fxp_functions_0_aadd_7_a62),
	.shareout());
defparam fxp_functions_0_aadd_7_a61.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a61.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a66(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a66_sumout),
	.cout(fxp_functions_0_aadd_7_a67),
	.shareout());
defparam fxp_functions_0_aadd_7_a66.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a66.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a71(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a14_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a71_sumout),
	.cout(fxp_functions_0_aadd_7_a72),
	.shareout());
defparam fxp_functions_0_aadd_7_a71.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a71.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a76(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a15_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a76_sumout),
	.cout(fxp_functions_0_aadd_7_a77),
	.shareout());
defparam fxp_functions_0_aadd_7_a76.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a76.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a81(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a16_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a81_sumout),
	.cout(fxp_functions_0_aadd_7_a82),
	.shareout());
defparam fxp_functions_0_aadd_7_a81.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a81.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a86(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a17_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a86_sumout),
	.cout(fxp_functions_0_aadd_7_a87),
	.shareout());
defparam fxp_functions_0_aadd_7_a86.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a86.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a91(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a18_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a91_sumout),
	.cout(fxp_functions_0_aadd_7_a92),
	.shareout());
defparam fxp_functions_0_aadd_7_a91.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a91.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a96(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a19_a),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a96_sumout),
	.cout(fxp_functions_0_aadd_7_a97),
	.shareout());
defparam fxp_functions_0_aadd_7_a96.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a96.lut_mask = 64'h00000000005555AA;
defparam fxp_functions_0_aadd_7_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a101(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a101_sumout),
	.cout(fxp_functions_0_aadd_7_a102),
	.shareout());
defparam fxp_functions_0_aadd_7_a101.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a101.lut_mask = 64'h0000000011116666;
defparam fxp_functions_0_aadd_7_a101.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_7_a106(
	.dataa(!fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq),
	.datab(!fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a20_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aadd_7_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aadd_7_a106_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_7_a106.extended_lut = "off";
defparam fxp_functions_0_aadd_7_a106.lut_mask = 64'h0000000000006666;
defparam fxp_functions_0_aadd_7_a106.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_1_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_9_a172(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aadd_9_a172_cout),
	.shareout());
defparam fxp_functions_0_aadd_9_a172.extended_lut = "off";
defparam fxp_functions_0_aadd_9_a172.lut_mask = 64'h00000000000F0FF0;
defparam fxp_functions_0_aadd_9_a172.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a12_a_a0_a.power_up = "dont_care";

fourteennm_mac fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0(
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.dfxlfsrena(vcc),
	.dfxmisrena(vcc),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a_aq}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a_aq,
fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a_aq,fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a_aq}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({clk,clk,clk}),
	.clr({rst,rst}),
	.ena({fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout,fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout}),
	.scanin(27'b000000000000000000000000000),
	.chainin(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.dftout(),
	.resulta(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0_RESULTA_bus),
	.resultb(),
	.scanout(),
	.chainout());
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.accum_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.accum_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.accumulate_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.ax_clock = "0";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.ax_width = 14;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.ay_scan_in_clock = "0";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.ay_scan_in_width = 14;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.ay_use_scan_in = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.az_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.bx_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.by_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.by_use_scan_in = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.bz_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.chainout_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.clear_type = "sclr";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_0 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_1 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_2 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_3 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_4 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_5 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_6 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_a_7 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_0 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_1 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_2 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_3 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_4 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_5 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_6 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_b_7 = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_sel_a_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.coef_sel_b_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.delay_scan_out_ay = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.delay_scan_out_by = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.enable_double_accum = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.input_pipeline_clock = "2";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.input_systolic_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.load_const_2nd_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.load_const_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.load_const_pipeline_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.load_const_value = 0;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.negate_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.operand_source_max = "input";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.operand_source_may = "input";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.operand_source_mbx = "input";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.operand_source_mby = "input";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.operation_mode = "m18x18_full";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.output_clock = "1";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.preadder_subtract_a = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.preadder_subtract_b = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.result_a_width = 28;
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.second_pipeline_clock = "2";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.signed_max = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.signed_may = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.signed_mbx = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.signed_mby = "false";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.sub_clock = "none";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_DSP0.use_chainadder = "false";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "9E020390CEC6182B9667F3A2C30A3E343FE385FF3A54CF98840D9131A6527CC7";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "B4BAA23432459D1DFF913D4EA55716A5E2F21B05765CA489C742459A7A22BAEB";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "63FA2D14F2E6A40201D02624C7E547EBFBFD2F90230C7B58E2AA2FB49C0B882A";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "E14787EBF3CC5C3F86846BC2B547C7EC1E0DC4D834C1306CD89E28F71D03B0FF";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "BEEAC6B04A5AD8AC6BE2A0B9F86BD2DE16EAA6F80F25F6AA88CEAD975EE4B0A8";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "94E702CD78BB30729BBF0EEEE23B4073823FFBC98ED82F5945FA5DEBD5E296ED";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "8DB401A98653F541AC6BE4E4EBECE1745F11112A46D8F9F4F09EE022D94B79F7";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "8392AACE01C95980654C1DB7194FD58D615F5F497CCFBA22DD5A6DAFB8159371";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "2ADB330FFFC734AAB6700392AD8FCCA980CA60DD826F93EB363233245A22549D";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "CCE3C3F0003F0C666D2AAADB31F03C64AA93803B548F894C0D5DEA2299416D09";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "5A56A9555555A94B49B3331C3E0003E399B6AAAD98F078DAA99FE68B18D58351";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "39CE6733333364D9249696B56AAAAAB52D24CCCE1F0007C664B54B33E7CCAA61";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "07C1E0F0F0F0E3C71C718E731999999364925A5AB555556B492673C3FFC3992B";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "003FE00FF00FE03F03F07E0F0787878F1C71C6398CCCCCD92492D6A9556AD24D";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_first_bit_number = 14;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_first_bit_number = 14;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a14.mem_init0 = "00001FFFF0001FFF000FFE00FF807F80FC0FC1F87C3C3C38E38E3198CCD9B6DB";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_first_bit_number = 15;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_first_bit_number = 15;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a15.mem_init0 = "000000000FFFFFFF000001FFFF80007FFC003FF803FC03F81F81F0783C3871C7";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_first_bit_number = 16;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_first_bit_number = 16;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a16.mem_init0 = "0000000000000000FFFFFFFFFF80000003FFFFF80003FFF8007FF007FC07F03F";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_first_bit_number = 17;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_first_bit_number = 17;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a17.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFF80000000000007FFFFFFF800000FFFFC000FFF";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_first_bit_number = 18;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_first_bit_number = 18;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a18.mem_init0 = "000000000000000000000000007FFFFFFFFFFFFFFFFFFFF80000000003FFFFFF";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_first_bit_number = 19;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_first_bit_number = 19;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a19.mem_init0 = "000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFF";

fourteennm_ram_block fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC2_uid80_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.logical_ram_name = "fxp_functions_0|memoryC2_uid80_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_first_bit_number = 20;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_a_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_first_bit_number = 20;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.port_b_logical_ram_width = 21;
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC2_uid80_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a20.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai2020_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.first_bit_number = 8;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama8";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama8.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.first_bit_number = 9;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama9";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama9.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.first_bit_number = 10;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama10";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama10.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.first_bit_number = 11;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama11";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama11.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.first_bit_number = 12;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama12";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama12.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.first_bit_number = 13;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama13";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama13.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.first_bit_number = 14;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama14";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama14.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.first_bit_number = 15;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama15";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama15.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.first_bit_number = 16;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama16";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama16.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.first_bit_number = 17;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama17";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama17.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.first_bit_number = 18;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama18";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama18.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.first_bit_number = 19;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama19";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama19.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.first_bit_number = 20;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama20";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama20.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.first_bit_number = 21;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama21";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama21.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.first_bit_number = 22;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama22";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama22.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a13_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_4_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist4_yaddr_uid19_divider_merged_bit_select_c_10_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 23;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a_aq));
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist1_yAddr_uid19_divider_merged_bit_select_b_14_inputreg0_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a22_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a14_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aq_a_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a_aq));
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_wire_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_adataout_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai2032_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai2032_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai2032_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a23_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a15_a_a0_a.power_up = "dont_care";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_first_bit_number = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_first_bit_number = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a0.mem_init0 = "56A567A7E28AF8C3AA2DA8DBD82D68E98AD3FFA6FAA6153F5112C50126481150";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_first_bit_number = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_first_bit_number = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a1.mem_init0 = "A40996F3C456F544D93AB483072882267F14115AED8C2EF23E3677785E6F9D53";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_first_bit_number = 2;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_first_bit_number = 2;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a2.mem_init0 = "922D1EA4DE56F6BCAA7FB4C86F5F8505F2CB39185F451814AA5911A94075E3D0";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_first_bit_number = 3;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_first_bit_number = 3;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a3.mem_init0 = "59137FC6A5B4A604893540CD97EC1F093CB0566C865E14B7FE2F62EA01862046";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_first_bit_number = 4;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_first_bit_number = 4;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a4.mem_init0 = "6161850CF9D73F1955A42610EA06D1446A94C137BE4097798FDB6FFC24B1D20E";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_first_bit_number = 5;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_first_bit_number = 5;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a5.mem_init0 = "7E81F80F01E8381E1E3A38E10C771989B3269A5AD4EABD6B66C71FFFC6DAA93E";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_first_bit_number = 6;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_first_bit_number = 6;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a6.mem_init0 = "7FFE000FFE003FE01FC03F01F0781E0E3C38E39CE773264DB495AAAAADB66701";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_first_bit_number = 7;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_first_bit_number = 7;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a7.mem_init0 = "7FFFFFF000003FFFE0003FFE007FE00FC03F03E0F87C3871C719CCCCC924B5AA";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_first_bit_number = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_first_bit_number = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a8.mem_init0 = "7FFFFFFFFFFFC00000003FFFFF80000FFFC003FF007FC07E07E1F0F0F1C739CC";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_first_bit_number = 9;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_first_bit_number = 9;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a9.mem_init0 = "800000000000000000003FFFFFFFFFF0000003FFFF80007FF801FF00FE07C1F0";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_first_bit_number = 10;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_first_bit_number = 10;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a10.mem_init0 = "FFFFFFFFFFFFFFFFFFFFC00000000000000003FFFFFFFF800001FFFF0007FE00";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_first_bit_number = 11;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_first_bit_number = 11;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a11.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000001FFFFFFF80000";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_first_bit_number = 12;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_first_bit_number = 12;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a12.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000";

fourteennm_ram_block fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13(
	.clk0(clk),
	.clk1(clk),
	.aclr(gnd),
	.sclr(rst),
	.ena0(en[0]),
	.ena1(en[0]),
	.portaaddrstall(gnd),
	.portaaddrstall2(gnd),
	.portare(vcc),
	.portawe(gnd),
	.eccencbypass(gnd),
	.portbaddrstall(gnd),
	.portbaddrstall2(gnd),
	.portbre(vcc),
	.portbwe(gnd),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portaaddr2(1'b0),
	.portabyteenamasks(1'b1),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.eccencparity(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aMux_72_a0_combout,fxp_functions_0_aMux_72_a32_sumout,fxp_functions_0_aMux_72_a27_sumout,fxp_functions_0_aMux_72_a22_sumout,fxp_functions_0_aMux_72_a17_sumout,fxp_functions_0_aMux_72_a12_sumout,
fxp_functions_0_aMux_72_a7_sumout,fxp_functions_0_aMux_72_a2_sumout}),
	.portbaddr2(1'b0),
	.portbbyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portadataout(),
	.portbdataout(fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_input_clock_enable = "ena0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk0_output_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_input_clock_enable = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.clk1_output_clock_enable = "ena1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_offset_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.data_interleave_width_in_bits = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_coherent_read = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_ecc_encoder_bypass = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.enable_force_to_zero = "false";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file = "../../altera_fxp_functions_191/synth/Fix_Div_altera_fxp_functions_191_fy4uury_memoryC3_uid83_invTabGen_lutmem.hex";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.init_file_layout = "port_a";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.logical_ram_name = "fxp_functions_0|memoryC3_uid83_invTabGen_lutmem_dmem|auto_generated|altera_syncram_impl1|ALTERA_SYNCRAM";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mixed_port_feed_through_mode = "dont_care";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.operation_mode = "dual_port";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clear = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_out_clock = "none";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_first_bit_number = 13;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_a_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_clock = "clock0";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_address_width = 8;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clear = "sclear";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_out_clock = "clock1";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_data_width = 1;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_address = 0;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_first_bit_number = 13;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_last_address = 255;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_depth = 256;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.port_b_logical_ram_width = 14;
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.ram_block_type = "M20K";
defparam fxp_functions_0_amemoryC3_uid83_invTabGen_lutmem_dmem_aauto_generated_aaltera_syncram_impl1_aram_block2a13.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a22_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.first_bit_number = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama0";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama0.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai4258_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a.power_up = "dont_care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.first_bit_number = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama1";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama1.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.first_bit_number = 2;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama2";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama2.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.first_bit_number = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama3";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama3.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.first_bit_number = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama4";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama4.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.first_bit_number = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama5";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama5.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.first_bit_number = 6;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama6";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama6.mixed_port_feed_through_mode = "dont care";

fourteennm_mlab_cell fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7(
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq}),
	.portaaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq}),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq,
fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq}),
	.portbdataout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7_PORTBDATAOUT_bus));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.address_width = 3;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.data_width = 1;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_address = 0;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.first_bit_number = 7;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.init_file = "none";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.last_address = 4;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_depth = 5;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_name = "fxp_functions_0|redist0_yaddr_uid19_divider_merged_bit_select_b_7_mem_dmem|auto_generated|altera_syncram_impl1|lutrama7";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.logical_ram_width = 8;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_alutrama7.mixed_port_feed_through_mode = "dont care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_5_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a24_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a16_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a76_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_11_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_93_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ai6615_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a_aq));
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a25_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a17_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai4270_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai4270_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai4270_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_95_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_94_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a26_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a18_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_12_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a27_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a19_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a(
	.clk(clk),
	.d(denominator[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a_aq));
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a28_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a20_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a29_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a_aq));
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a21_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a30_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_anormYIsOne_uid16_divider_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a31_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_64_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a12_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a7_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a2_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a27_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a32_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a22_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a17_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a_aq));
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a_aq));
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a32_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_areduce_nor_18_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_ayIsZero_uid17_divider_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_1_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(rst),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a_aq));
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_delay_0_a31_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aMux_99_a2(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_99_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_99_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_99_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_99_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_99_a6(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_99_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_99_a6_sumout),
	.cout(fxp_functions_0_aMux_99_a7),
	.shareout());
defparam fxp_functions_0_aMux_99_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_99_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_99_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_100_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_99_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_100_a1_sumout),
	.cout(fxp_functions_0_aMux_100_a2),
	.shareout());
defparam fxp_functions_0_aMux_100_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_100_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_100_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_101_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a61_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_100_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_101_a1_sumout),
	.cout(fxp_functions_0_aMux_101_a2),
	.shareout());
defparam fxp_functions_0_aMux_101_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_101_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_101_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_102_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a60_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_101_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_102_a1_sumout),
	.cout(fxp_functions_0_aMux_102_a2),
	.shareout());
defparam fxp_functions_0_aMux_102_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_102_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_102_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_103_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a59_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_102_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_103_a1_sumout),
	.cout(fxp_functions_0_aMux_103_a2),
	.shareout());
defparam fxp_functions_0_aMux_103_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_103_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_103_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_104_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a58_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_103_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_104_a1_sumout),
	.cout(fxp_functions_0_aMux_104_a2),
	.shareout());
defparam fxp_functions_0_aMux_104_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_104_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_104_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_105_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a57_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_104_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_105_a1_sumout),
	.cout(fxp_functions_0_aMux_105_a2),
	.shareout());
defparam fxp_functions_0_aMux_105_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_105_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_105_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_106_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a56_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_105_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_106_a1_sumout),
	.cout(fxp_functions_0_aMux_106_a2),
	.shareout());
defparam fxp_functions_0_aMux_106_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_106_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_106_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_107_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a55_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_106_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_107_a1_sumout),
	.cout(fxp_functions_0_aMux_107_a2),
	.shareout());
defparam fxp_functions_0_aMux_107_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_107_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_107_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_108_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a54_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_107_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_108_a1_sumout),
	.cout(fxp_functions_0_aMux_108_a2),
	.shareout());
defparam fxp_functions_0_aMux_108_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_108_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_108_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_109_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a53_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_108_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_109_a1_sumout),
	.cout(fxp_functions_0_aMux_109_a2),
	.shareout());
defparam fxp_functions_0_aMux_109_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_109_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_109_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_110_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a52_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_109_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_110_a1_sumout),
	.cout(fxp_functions_0_aMux_110_a2),
	.shareout());
defparam fxp_functions_0_aMux_110_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_110_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_110_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_111_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a51_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_110_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_111_a1_sumout),
	.cout(fxp_functions_0_aMux_111_a2),
	.shareout());
defparam fxp_functions_0_aMux_111_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_111_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_111_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_112_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a50_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_111_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_112_a1_sumout),
	.cout(fxp_functions_0_aMux_112_a2),
	.shareout());
defparam fxp_functions_0_aMux_112_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_112_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_112_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_113_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a49_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_112_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_113_a1_sumout),
	.cout(fxp_functions_0_aMux_113_a2),
	.shareout());
defparam fxp_functions_0_aMux_113_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_113_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_113_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_114_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a48_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_113_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_114_a1_sumout),
	.cout(fxp_functions_0_aMux_114_a2),
	.shareout());
defparam fxp_functions_0_aMux_114_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_114_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_114_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_115_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a47_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_114_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_115_a1_sumout),
	.cout(fxp_functions_0_aMux_115_a2),
	.shareout());
defparam fxp_functions_0_aMux_115_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_115_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_115_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_116_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a46_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_115_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_116_a1_sumout),
	.cout(fxp_functions_0_aMux_116_a2),
	.shareout());
defparam fxp_functions_0_aMux_116_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_116_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_116_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_117_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_116_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_117_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_117_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_117_a1.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_117_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_118_a2(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a45_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_118_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_118_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_118_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_118_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_118_a6(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a44_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_118_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_118_a6_sumout),
	.cout(fxp_functions_0_aMux_118_a7),
	.shareout());
defparam fxp_functions_0_aMux_118_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_118_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_118_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_119_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a43_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_118_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_119_a1_sumout),
	.cout(fxp_functions_0_aMux_119_a2),
	.shareout());
defparam fxp_functions_0_aMux_119_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_119_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_119_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_120_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a42_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_119_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_120_a1_sumout),
	.cout(fxp_functions_0_aMux_120_a2),
	.shareout());
defparam fxp_functions_0_aMux_120_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_120_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_120_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_121_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a41_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_120_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_121_a1_sumout),
	.cout(fxp_functions_0_aMux_121_a2),
	.shareout());
defparam fxp_functions_0_aMux_121_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_121_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_121_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_122_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a40_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_121_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_122_a1_sumout),
	.cout(fxp_functions_0_aMux_122_a2),
	.shareout());
defparam fxp_functions_0_aMux_122_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_122_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_122_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_123_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a39_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_122_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_123_a1_sumout),
	.cout(fxp_functions_0_aMux_123_a2),
	.shareout());
defparam fxp_functions_0_aMux_123_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_123_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_123_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_124_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a38_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_123_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_124_a1_sumout),
	.cout(fxp_functions_0_aMux_124_a2),
	.shareout());
defparam fxp_functions_0_aMux_124_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_124_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_124_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_125_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a37_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_124_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_125_a1_sumout),
	.cout(fxp_functions_0_aMux_125_a2),
	.shareout());
defparam fxp_functions_0_aMux_125_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_125_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_125_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a13(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a36_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_125_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai8489_a13_sumout),
	.cout(fxp_functions_0_ai8489_a14),
	.shareout());
defparam fxp_functions_0_ai8489_a13.extended_lut = "off";
defparam fxp_functions_0_ai8489_a13.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai8489_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a18(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a35_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai8489_a14),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai8489_a18_sumout),
	.cout(fxp_functions_0_ai8489_a19),
	.shareout());
defparam fxp_functions_0_ai8489_a18.extended_lut = "off";
defparam fxp_functions_0_ai8489_a18.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai8489_a18.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a23(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a32_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a34_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai8489_a19),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai8489_a23_sumout),
	.cout(fxp_functions_0_ai8489_a24),
	.shareout());
defparam fxp_functions_0_ai8489_a23.extended_lut = "off";
defparam fxp_functions_0_ai8489_a23.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai8489_a23.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a28(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a31_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a33_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai8489_a24),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai8489_a28_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a28.extended_lut = "off";
defparam fxp_functions_0_ai8489_a28.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_ai8489_a28.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_48_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_20_a0_combout),
	.datad(!fxp_functions_0_aMux_28_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_48_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_48_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_48_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_48_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_48_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_16_a0_combout),
	.datad(!fxp_functions_0_aMux_24_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_48_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_48_a6_sumout),
	.cout(fxp_functions_0_aMux_48_a7),
	.shareout());
defparam fxp_functions_0_aMux_48_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_48_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_48_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_44_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_12_a1_combout),
	.datad(!fxp_functions_0_aMux_20_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_48_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_44_a1_sumout),
	.cout(fxp_functions_0_aMux_44_a2),
	.shareout());
defparam fxp_functions_0_aMux_44_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_44_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_44_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a19(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_8_a1_combout),
	.datad(!fxp_functions_0_aMux_16_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_44_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_40_a19_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a19.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a19.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_40_a19.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_50_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_22_a0_combout),
	.datad(!fxp_functions_0_aMux_30_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_50_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_50_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_50_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_50_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_50_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_18_a0_combout),
	.datad(!fxp_functions_0_aMux_26_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_50_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_50_a6_sumout),
	.cout(fxp_functions_0_aMux_50_a7),
	.shareout());
defparam fxp_functions_0_aMux_50_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_50_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_50_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_46_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_14_a1_combout),
	.datad(!fxp_functions_0_aMux_22_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_50_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_46_a1_sumout),
	.cout(fxp_functions_0_aMux_46_a2),
	.shareout());
defparam fxp_functions_0_aMux_46_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_46_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_46_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_42_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_10_a1_combout),
	.datad(!fxp_functions_0_aMux_18_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_46_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_42_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_42_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_42_a1.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_42_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_49_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_21_a0_combout),
	.datad(!fxp_functions_0_aMux_29_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_49_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_49_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_49_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_49_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_49_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_17_a0_combout),
	.datad(!fxp_functions_0_aMux_25_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_49_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_49_a6_sumout),
	.cout(fxp_functions_0_aMux_49_a7),
	.shareout());
defparam fxp_functions_0_aMux_49_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_49_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_49_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_45_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_13_a1_combout),
	.datad(!fxp_functions_0_aMux_21_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_49_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_45_a1_sumout),
	.cout(fxp_functions_0_aMux_45_a2),
	.shareout());
defparam fxp_functions_0_aMux_45_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_45_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_45_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_41_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_9_a1_combout),
	.datad(!fxp_functions_0_aMux_17_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_45_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_41_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_41_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_41_a1.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_41_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_51_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_23_a0_combout),
	.datad(!fxp_functions_0_aMux_31_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_aMux_51_a2_cout),
	.shareout());
defparam fxp_functions_0_aMux_51_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_51_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_aMux_51_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_51_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_19_a0_combout),
	.datad(!fxp_functions_0_aMux_27_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_51_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_51_a6_sumout),
	.cout(fxp_functions_0_aMux_51_a7),
	.shareout());
defparam fxp_functions_0_aMux_51_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_51_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_51_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_47_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_15_a1_combout),
	.datad(!fxp_functions_0_aMux_23_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_51_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_47_a1_sumout),
	.cout(fxp_functions_0_aMux_47_a2),
	.shareout());
defparam fxp_functions_0_aMux_47_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_47_a1.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_47_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_43_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aMux_11_a1_combout),
	.datad(!fxp_functions_0_aMux_19_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_47_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_43_a1_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_43_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_43_a1.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_43_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_61_a0_combout),
	.datad(!fxp_functions_0_aMux_63_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_ai6615_a2_cout),
	.shareout());
defparam fxp_functions_0_ai6615_a2.extended_lut = "off";
defparam fxp_functions_0_ai6615_a2.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_ai6615_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_60_a0_combout),
	.datad(!fxp_functions_0_aMux_62_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a2_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a6_sumout),
	.cout(fxp_functions_0_ai6615_a7),
	.shareout());
defparam fxp_functions_0_ai6615_a6.extended_lut = "off";
defparam fxp_functions_0_ai6615_a6.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a11(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_59_a1_combout),
	.datad(!fxp_functions_0_aMux_61_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a11_sumout),
	.cout(fxp_functions_0_ai6615_a12),
	.shareout());
defparam fxp_functions_0_ai6615_a11.extended_lut = "off";
defparam fxp_functions_0_ai6615_a11.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a16(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_58_a1_combout),
	.datad(!fxp_functions_0_aMux_60_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a16_sumout),
	.cout(fxp_functions_0_ai6615_a17),
	.shareout());
defparam fxp_functions_0_ai6615_a16.extended_lut = "off";
defparam fxp_functions_0_ai6615_a16.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a21(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_57_a1_combout),
	.datad(!fxp_functions_0_aMux_59_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a21_sumout),
	.cout(fxp_functions_0_ai6615_a22),
	.shareout());
defparam fxp_functions_0_ai6615_a21.extended_lut = "off";
defparam fxp_functions_0_ai6615_a21.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a26(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_56_a1_combout),
	.datad(!fxp_functions_0_aMux_58_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a26_sumout),
	.cout(fxp_functions_0_ai6615_a27),
	.shareout());
defparam fxp_functions_0_ai6615_a26.extended_lut = "off";
defparam fxp_functions_0_ai6615_a26.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a31(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_55_a0_combout),
	.datad(!fxp_functions_0_aMux_57_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a31_sumout),
	.cout(fxp_functions_0_ai6615_a32),
	.shareout());
defparam fxp_functions_0_ai6615_a31.extended_lut = "off";
defparam fxp_functions_0_ai6615_a31.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a36(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_54_a0_combout),
	.datad(!fxp_functions_0_aMux_56_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a36_sumout),
	.cout(fxp_functions_0_ai6615_a37),
	.shareout());
defparam fxp_functions_0_ai6615_a36.extended_lut = "off";
defparam fxp_functions_0_ai6615_a36.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a36.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a41(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_53_a0_combout),
	.datad(!fxp_functions_0_aMux_55_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a41_sumout),
	.cout(fxp_functions_0_ai6615_a42),
	.shareout());
defparam fxp_functions_0_ai6615_a41.extended_lut = "off";
defparam fxp_functions_0_ai6615_a41.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a41.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a46(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_52_a0_combout),
	.datad(!fxp_functions_0_aMux_54_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a46_sumout),
	.cout(fxp_functions_0_ai6615_a47),
	.shareout());
defparam fxp_functions_0_ai6615_a46.extended_lut = "off";
defparam fxp_functions_0_ai6615_a46.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a46.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a51(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_51_a6_sumout),
	.datad(!fxp_functions_0_aMux_53_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a51_sumout),
	.cout(fxp_functions_0_ai6615_a52),
	.shareout());
defparam fxp_functions_0_ai6615_a51.extended_lut = "off";
defparam fxp_functions_0_ai6615_a51.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a51.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a56(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_50_a6_sumout),
	.datad(!fxp_functions_0_aMux_52_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a56_sumout),
	.cout(fxp_functions_0_ai6615_a57),
	.shareout());
defparam fxp_functions_0_ai6615_a56.extended_lut = "off";
defparam fxp_functions_0_ai6615_a56.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a56.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a61(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_49_a6_sumout),
	.datad(!fxp_functions_0_aMux_51_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a61_sumout),
	.cout(fxp_functions_0_ai6615_a62),
	.shareout());
defparam fxp_functions_0_ai6615_a61.extended_lut = "off";
defparam fxp_functions_0_ai6615_a61.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a61.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a66(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_48_a6_sumout),
	.datad(!fxp_functions_0_aMux_50_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a66_sumout),
	.cout(fxp_functions_0_ai6615_a67),
	.shareout());
defparam fxp_functions_0_ai6615_a66.extended_lut = "off";
defparam fxp_functions_0_ai6615_a66.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a66.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a71(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_47_a1_sumout),
	.datad(!fxp_functions_0_aMux_49_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a71_sumout),
	.cout(fxp_functions_0_ai6615_a72),
	.shareout());
defparam fxp_functions_0_ai6615_a71.extended_lut = "off";
defparam fxp_functions_0_ai6615_a71.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a71.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a76(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_46_a1_sumout),
	.datad(!fxp_functions_0_aMux_48_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a76_sumout),
	.cout(fxp_functions_0_ai6615_a77),
	.shareout());
defparam fxp_functions_0_ai6615_a76.extended_lut = "off";
defparam fxp_functions_0_ai6615_a76.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a76.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a81(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_45_a1_sumout),
	.datad(!fxp_functions_0_aMux_47_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a81_sumout),
	.cout(fxp_functions_0_ai6615_a82),
	.shareout());
defparam fxp_functions_0_ai6615_a81.extended_lut = "off";
defparam fxp_functions_0_ai6615_a81.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a81.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a86(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_44_a1_sumout),
	.datad(!fxp_functions_0_aMux_46_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a86_sumout),
	.cout(fxp_functions_0_ai6615_a87),
	.shareout());
defparam fxp_functions_0_ai6615_a86.extended_lut = "off";
defparam fxp_functions_0_ai6615_a86.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a86.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a91(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_43_a1_sumout),
	.datad(!fxp_functions_0_aMux_45_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a91_sumout),
	.cout(fxp_functions_0_ai6615_a92),
	.shareout());
defparam fxp_functions_0_ai6615_a91.extended_lut = "off";
defparam fxp_functions_0_ai6615_a91.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a91.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a96(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_42_a1_sumout),
	.datad(!fxp_functions_0_aMux_44_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a96_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6615_a96.extended_lut = "off";
defparam fxp_functions_0_ai6615_a96.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_ai6615_a96.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a102(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_42_a1_sumout),
	.datad(!fxp_functions_0_aMux_44_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fxp_functions_0_ai6615_a102_cout),
	.shareout());
defparam fxp_functions_0_ai6615_a102.extended_lut = "off";
defparam fxp_functions_0_ai6615_a102.lut_mask = 64'h0000000004150000;
defparam fxp_functions_0_ai6615_a102.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6615_a106(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_41_a1_sumout),
	.datad(!fxp_functions_0_aMux_43_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a102_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_ai6615_a106_sumout),
	.cout(fxp_functions_0_ai6615_a107),
	.shareout());
defparam fxp_functions_0_ai6615_a106.extended_lut = "off";
defparam fxp_functions_0_ai6615_a106.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_ai6615_a106.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a19_sumout),
	.datad(!fxp_functions_0_aMux_42_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_ai6615_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a2_sumout),
	.cout(fxp_functions_0_aMux_72_a3),
	.shareout());
defparam fxp_functions_0_aMux_72_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a2.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a7(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a2_combout),
	.datad(!fxp_functions_0_aMux_41_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a3),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a7_sumout),
	.cout(fxp_functions_0_aMux_72_a8),
	.shareout());
defparam fxp_functions_0_aMux_72_a7.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a7.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a12(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a5_combout),
	.datad(!fxp_functions_0_aMux_40_a19_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a8),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a12_sumout),
	.cout(fxp_functions_0_aMux_72_a13),
	.shareout());
defparam fxp_functions_0_aMux_72_a12.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a12.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a17(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a8_combout),
	.datad(!fxp_functions_0_aMux_40_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a13),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a17_sumout),
	.cout(fxp_functions_0_aMux_72_a18),
	.shareout());
defparam fxp_functions_0_aMux_72_a17.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a17.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a22(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a9_combout),
	.datad(!fxp_functions_0_aMux_40_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a18),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a22_sumout),
	.cout(fxp_functions_0_aMux_72_a23),
	.shareout());
defparam fxp_functions_0_aMux_72_a22.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a22.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a27(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a12_combout),
	.datad(!fxp_functions_0_aMux_40_a8_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a23),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a27_sumout),
	.cout(fxp_functions_0_aMux_72_a28),
	.shareout());
defparam fxp_functions_0_aMux_72_a27.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a27.lut_mask = 64'h000000000415082A;
defparam fxp_functions_0_aMux_72_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a32(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aMux_40_a14_combout),
	.datad(!fxp_functions_0_aMux_40_a9_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fxp_functions_0_aMux_72_a28),
	.sharein(gnd),
	.combout(),
	.sumout(fxp_functions_0_aMux_72_a32_sumout),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_72_a32.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a32.lut_mask = 64'h000000000000082A;
defparam fxp_functions_0_aMux_72_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_64_a1(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_40_a13_combout),
	.datad(!fxp_functions_0_aMux_40_a10_combout),
	.datae(!fxp_functions_0_aMux_40_a17_combout),
	.dataf(!fxp_functions_0_aMux_32_a2_combout),
	.datag(!fxp_functions_0_aMux_32_a3_combout),
	.datah(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_64_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_64_a1.extended_lut = "on";
defparam fxp_functions_0_aMux_64_a1.lut_mask = 64'h03CF03CF0C4C3F7F;
defparam fxp_functions_0_aMux_64_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_32_a3(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a_aq),
	.datae(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.dataf(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datag(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a_aq),
	.datah(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_32_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_32_a3.extended_lut = "on";
defparam fxp_functions_0_aMux_32_a3.lut_mask = 64'h05F5000003F30000;
defparam fxp_functions_0_aMux_32_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_64_a6(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_40_a11_combout),
	.datad(!fxp_functions_0_aMux_40_a10_combout),
	.datae(!fxp_functions_0_aMux_40_a16_combout),
	.dataf(!fxp_functions_0_aMux_40_a15_combout),
	.datag(!fxp_functions_0_aMux_40_a23_combout),
	.datah(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_64_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_64_a6.extended_lut = "on";
defparam fxp_functions_0_aMux_64_a6.lut_mask = 64'h03CF03CF0C4C3F7F;
defparam fxp_functions_0_aMux_64_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a23(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a_aq),
	.datae(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.dataf(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datag(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a_aq),
	.datah(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a23.extended_lut = "on";
defparam fxp_functions_0_aMux_40_a23.lut_mask = 64'h05F5000003F30000;
defparam fxp_functions_0_aMux_40_a23.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a34(
	.dataa(!fxp_functions_0_aMux_98_a0_combout),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datac(!fxp_functions_0_aMux_102_a1_sumout),
	.datad(!fxp_functions_0_aMux_110_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_106_a1_sumout),
	.datag(!fxp_functions_0_aMux_114_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a34_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a34.extended_lut = "on";
defparam fxp_functions_0_ai8489_a34.lut_mask = 64'h03CF444403CF0000;
defparam fxp_functions_0_ai8489_a34.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a39(
	.dataa(!fxp_functions_0_aMux_99_a6_sumout),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datac(!fxp_functions_0_aMux_103_a1_sumout),
	.datad(!fxp_functions_0_aMux_111_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_107_a1_sumout),
	.datag(!fxp_functions_0_aMux_115_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a39_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a39.extended_lut = "on";
defparam fxp_functions_0_ai8489_a39.lut_mask = 64'h03CF444403CF0000;
defparam fxp_functions_0_ai8489_a39.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a44(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_167_a1_combout),
	.datac(!fxp_functions_0_aMux_106_a1_sumout),
	.datad(!fxp_functions_0_aMux_114_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_110_a1_sumout),
	.datag(!fxp_functions_0_aMux_118_a6_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a44_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a44.extended_lut = "on";
defparam fxp_functions_0_ai8489_a44.lut_mask = 64'h05AF333305AF3333;
defparam fxp_functions_0_ai8489_a44.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a49(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_168_a1_combout),
	.datac(!fxp_functions_0_aMux_107_a1_sumout),
	.datad(!fxp_functions_0_aMux_115_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_111_a1_sumout),
	.datag(!fxp_functions_0_aMux_119_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a49_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a49.extended_lut = "on";
defparam fxp_functions_0_ai8489_a49.lut_mask = 64'h05AF333305AF3333;
defparam fxp_functions_0_ai8489_a49.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a54(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datab(!fxp_functions_0_aMux_169_a0_combout),
	.datac(!fxp_functions_0_aMux_112_a1_sumout),
	.datad(!fxp_functions_0_aMux_108_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_120_a1_sumout),
	.datag(!fxp_functions_0_aMux_116_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a54_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a54.extended_lut = "on";
defparam fxp_functions_0_ai8489_a54.lut_mask = 64'h0A5F33330A5F3333;
defparam fxp_functions_0_ai8489_a54.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a59(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datab(!fxp_functions_0_aMux_170_a0_combout),
	.datac(!fxp_functions_0_aMux_113_a1_sumout),
	.datad(!fxp_functions_0_aMux_109_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_121_a1_sumout),
	.datag(!fxp_functions_0_aMux_117_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a59_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a59.extended_lut = "on";
defparam fxp_functions_0_ai8489_a59.lut_mask = 64'h0A5F33330A5F3333;
defparam fxp_functions_0_ai8489_a59.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a64(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_171_a0_combout),
	.datac(!fxp_functions_0_aMux_110_a1_sumout),
	.datad(!fxp_functions_0_aMux_118_a6_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_122_a1_sumout),
	.datag(!fxp_functions_0_aMux_114_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a64_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a64.extended_lut = "on";
defparam fxp_functions_0_ai8489_a64.lut_mask = 64'h0A5F333305AF3333;
defparam fxp_functions_0_ai8489_a64.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a69(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_172_a0_combout),
	.datac(!fxp_functions_0_aMux_111_a1_sumout),
	.datad(!fxp_functions_0_aMux_119_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_123_a1_sumout),
	.datag(!fxp_functions_0_aMux_115_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a69_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a69.extended_lut = "on";
defparam fxp_functions_0_ai8489_a69.lut_mask = 64'h0A5F333305AF3333;
defparam fxp_functions_0_ai8489_a69.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a74(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_173_a0_combout),
	.datac(!fxp_functions_0_aMux_120_a1_sumout),
	.datad(!fxp_functions_0_aMux_112_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_124_a1_sumout),
	.datag(!fxp_functions_0_aMux_116_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a74_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a74.extended_lut = "on";
defparam fxp_functions_0_ai8489_a74.lut_mask = 64'h0A5F33330A5F3333;
defparam fxp_functions_0_ai8489_a74.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a79(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_aMux_174_a0_combout),
	.datac(!fxp_functions_0_aMux_121_a1_sumout),
	.datad(!fxp_functions_0_aMux_113_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.dataf(!fxp_functions_0_aMux_125_a1_sumout),
	.datag(!fxp_functions_0_aMux_117_a1_sumout),
	.datah(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a79_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a79.extended_lut = "on";
defparam fxp_functions_0_ai8489_a79.lut_mask = 64'h0A5F33330A5F3333;
defparam fxp_functions_0_ai8489_a79.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0(
	.dataa(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a3_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a4_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a5_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a6_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a7_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a8_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a9_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a10_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a11_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a12_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a13_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a14_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a15_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a16_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a17_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a18_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a19_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a20_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a21_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a22_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a23_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a24_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a25_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a26_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a27_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a28_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a29_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a30_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31(
	.dataa(!fxp_functions_0_aredist17_yIsZero_uid17_divider_q_34_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist15_prodPostRightShiftPostRndRange_uid35_divider_b_1_q_a31_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31.extended_lut = "off";
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0.extended_lut = "off";
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aMux_177_a0(
	.dataa(!fxp_functions_0_aMux_112_a1_sumout),
	.datab(!fxp_functions_0_aMux_104_a1_sumout),
	.datac(!fxp_functions_0_aMux_108_a1_sumout),
	.datad(!fxp_functions_0_aMux_100_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_177_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_177_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_177_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_177_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a0(
	.dataa(!fxp_functions_0_ai8489_a23_sumout),
	.datab(!fxp_functions_0_aMux_120_a1_sumout),
	.datac(!fxp_functions_0_aMux_124_a1_sumout),
	.datad(!fxp_functions_0_aMux_116_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a0.extended_lut = "off";
defparam fxp_functions_0_ai8489_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_ai8489_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a1(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datad(!fxp_functions_0_aMux_177_a0_combout),
	.datae(!fxp_functions_0_ai8489_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a1.extended_lut = "off";
defparam fxp_functions_0_ai8489_a1.lut_mask = 64'h002080A0002080A0;
defparam fxp_functions_0_ai8489_a1.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai8489_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a_aq));
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a0(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a14_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a11_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a0.lut_mask = 64'h0101010101010101;
defparam fxp_functions_0_areduce_nor_0_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a1(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a10_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a9_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a7_a_aq),
	.datae(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a5_a_aq),
	.dataf(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a6_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a1.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a1.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_0_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a2(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a13_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a32_a_aq),
	.datae(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a30_a_aq),
	.dataf(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a31_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a2.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a2.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_0_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a3(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a29_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a28_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a27_a_aq),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a26_a_aq),
	.datae(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a24_a_aq),
	.dataf(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a25_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a3.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a3.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_0_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a4(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a17_a_aq),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a16_a_aq),
	.datae(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_aq),
	.dataf(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a4.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a4.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_0_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0_a5(
	.dataa(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a23_a_aq),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a22_a_aq),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a21_a_aq),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a20_a_aq),
	.datae(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a18_a_aq),
	.dataf(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a19_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0_a5.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0_a5.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_0_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_0(
	.dataa(!fxp_functions_0_areduce_nor_0_a0_combout),
	.datab(!fxp_functions_0_areduce_nor_0_a1_combout),
	.datac(!fxp_functions_0_areduce_nor_0_a2_combout),
	.datad(!fxp_functions_0_areduce_nor_0_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_0_a4_combout),
	.dataf(!fxp_functions_0_areduce_nor_0_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_0_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_0.lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam fxp_functions_0_areduce_nor_0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_176_a0(
	.dataa(!fxp_functions_0_aMux_111_a1_sumout),
	.datab(!fxp_functions_0_aMux_103_a1_sumout),
	.datac(!fxp_functions_0_aMux_107_a1_sumout),
	.datad(!fxp_functions_0_aMux_99_a6_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_176_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_176_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_176_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_176_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datad(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0.lut_mask = 64'h08AA000008AA0000;
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datad(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1.lut_mask = 64'hA2AA0000A2AA0000;
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a2(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_115_a1_sumout),
	.datad(!fxp_functions_0_aMux_119_a1_sumout),
	.datae(!fxp_functions_0_ai8489_a18_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a2.extended_lut = "off";
defparam fxp_functions_0_ai8489_a2.lut_mask = 64'h03478BCF03478BCF;
defparam fxp_functions_0_ai8489_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a3(
	.dataa(!fxp_functions_0_aMux_123_a1_sumout),
	.datab(!fxp_functions_0_aMux_176_a0_combout),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0_combout),
	.datad(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1_combout),
	.datae(!fxp_functions_0_ai8489_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a3.extended_lut = "off";
defparam fxp_functions_0_ai8489_a3.lut_mask = 64'h050305F3050305F3;
defparam fxp_functions_0_ai8489_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a4(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_114_a1_sumout),
	.datad(!fxp_functions_0_aMux_118_a6_sumout),
	.datae(!fxp_functions_0_ai8489_a13_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a4.extended_lut = "off";
defparam fxp_functions_0_ai8489_a4.lut_mask = 64'h03478BCF03478BCF;
defparam fxp_functions_0_ai8489_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_98_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a62_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq),
	.datae(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_98_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_98_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_98_a0.lut_mask = 64'h082A4C6E082A4C6E;
defparam fxp_functions_0_aMux_98_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_175_a0(
	.dataa(!fxp_functions_0_aMux_110_a1_sumout),
	.datab(!fxp_functions_0_aMux_102_a1_sumout),
	.datac(!fxp_functions_0_aMux_106_a1_sumout),
	.datad(!fxp_functions_0_aMux_98_a0_combout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_175_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_175_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_175_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_175_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a5(
	.dataa(!fxp_functions_0_aMux_122_a1_sumout),
	.datab(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a0_combout),
	.datac(!fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a3_a_a1_combout),
	.datad(!fxp_functions_0_ai8489_a4_combout),
	.datae(!fxp_functions_0_aMux_175_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a5.extended_lut = "off";
defparam fxp_functions_0_ai8489_a5.lut_mask = 64'h101C131F101C131F;
defparam fxp_functions_0_ai8489_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_97_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq),
	.datad(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_97_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_97_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_97_a1.lut_mask = 64'h082A082A082A082A;
defparam fxp_functions_0_aMux_97_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_174_a0(
	.dataa(!fxp_functions_0_aMux_109_a1_sumout),
	.datab(!fxp_functions_0_aMux_101_a1_sumout),
	.datac(!fxp_functions_0_aMux_105_a1_sumout),
	.datad(!fxp_functions_0_aMux_97_a1_combout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_174_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_174_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_174_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_174_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_96_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_96_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_96_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_96_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_96_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_173_a0(
	.dataa(!fxp_functions_0_aMux_108_a1_sumout),
	.datab(!fxp_functions_0_aMux_100_a1_sumout),
	.datac(!fxp_functions_0_aMux_104_a1_sumout),
	.datad(!fxp_functions_0_aMux_96_a0_combout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_173_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_173_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_173_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_173_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_172_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_103_a1_sumout),
	.datad(!fxp_functions_0_aMux_107_a1_sumout),
	.datae(!fxp_functions_0_aMux_99_a6_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_172_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_172_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_172_a0.lut_mask = 64'h028A46CE028A46CE;
defparam fxp_functions_0_aMux_172_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_171_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_102_a1_sumout),
	.datad(!fxp_functions_0_aMux_106_a1_sumout),
	.datae(!fxp_functions_0_aMux_98_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_171_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_171_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_171_a0.lut_mask = 64'h028A46CE028A46CE;
defparam fxp_functions_0_aMux_171_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_170_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_101_a1_sumout),
	.datad(!fxp_functions_0_aMux_105_a1_sumout),
	.datae(!fxp_functions_0_aMux_97_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_170_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_170_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_170_a0.lut_mask = 64'h028A46CE028A46CE;
defparam fxp_functions_0_aMux_170_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_169_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_104_a1_sumout),
	.datad(!fxp_functions_0_aMux_100_a1_sumout),
	.datae(!fxp_functions_0_aMux_96_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_169_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_169_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_169_a0.lut_mask = 64'h082A4C6E082A4C6E;
defparam fxp_functions_0_aMux_169_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_168_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_103_a1_sumout),
	.datad(!fxp_functions_0_aMux_99_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_168_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_168_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_168_a1.lut_mask = 64'h082A082A082A082A;
defparam fxp_functions_0_aMux_168_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_167_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_102_a1_sumout),
	.datad(!fxp_functions_0_aMux_98_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_167_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_167_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_167_a1.lut_mask = 64'h082A082A082A082A;
defparam fxp_functions_0_aMux_167_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_166_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_101_a1_sumout),
	.datad(!fxp_functions_0_aMux_97_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_166_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_166_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_166_a1.lut_mask = 64'h082A082A082A082A;
defparam fxp_functions_0_aMux_166_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a6(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datab(!fxp_functions_0_aMux_166_a1_combout),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datad(!fxp_functions_0_aMux_113_a1_sumout),
	.datae(!fxp_functions_0_aMux_117_a1_sumout),
	.dataf(!fxp_functions_0_ai8489_a32_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a6.extended_lut = "off";
defparam fxp_functions_0_ai8489_a6.lut_mask = 64'h11B111B11B1BBBBB;
defparam fxp_functions_0_ai8489_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_165_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_100_a1_sumout),
	.datad(!fxp_functions_0_aMux_96_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_165_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_165_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_165_a1.lut_mask = 64'h082A082A082A082A;
defparam fxp_functions_0_aMux_165_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a7(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datab(!fxp_functions_0_aMux_165_a1_combout),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datad(!fxp_functions_0_aMux_112_a1_sumout),
	.datae(!fxp_functions_0_aMux_116_a1_sumout),
	.dataf(!fxp_functions_0_ai8489_a33_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a7.extended_lut = "off";
defparam fxp_functions_0_ai8489_a7.lut_mask = 64'h11B111B11B1BBBBB;
defparam fxp_functions_0_ai8489_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_162_a0(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_162_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_162_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_162_a0.lut_mask = 64'h8888888888888888;
defparam fxp_functions_0_aMux_162_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_164_a0(
	.dataa(!fxp_functions_0_aMux_99_a6_sumout),
	.datab(!fxp_functions_0_aMux_162_a0_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_164_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_164_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_164_a0.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aMux_164_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_163_a0(
	.dataa(!fxp_functions_0_aMux_162_a0_combout),
	.datab(!fxp_functions_0_aMux_98_a0_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_163_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_163_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_163_a0.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aMux_163_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_178_a0(
	.dataa(!fxp_functions_0_aMux_113_a1_sumout),
	.datab(!fxp_functions_0_aMux_105_a1_sumout),
	.datac(!fxp_functions_0_aMux_109_a1_sumout),
	.datad(!fxp_functions_0_aMux_101_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_178_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_178_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_178_a0.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_aMux_178_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_162_a1(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a1_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a0_a_aq),
	.datac(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a63_a_aq),
	.datad(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.dataf(!fxp_functions_0_aprodXInvY_uid27_divider_sums_result_add_0_0_o_a64_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_162_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_162_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_162_a1.lut_mask = 64'h080000002A000000;
defparam fxp_functions_0_aMux_162_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a8(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datad(!fxp_functions_0_aMux_178_a0_combout),
	.datae(!fxp_functions_0_aMux_162_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a8.extended_lut = "off";
defparam fxp_functions_0_ai8489_a8.lut_mask = 64'h008020A0008020A0;
defparam fxp_functions_0_ai8489_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a9(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datad(!fxp_functions_0_aMux_162_a0_combout),
	.datae(!fxp_functions_0_aMux_177_a0_combout),
	.dataf(!fxp_functions_0_aMux_96_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a9.extended_lut = "off";
defparam fxp_functions_0_ai8489_a9.lut_mask = 64'h00008080002080A0;
defparam fxp_functions_0_ai8489_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3.extended_lut = "off";
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam fxp_functions_0_aredist16_prodPostRightShiftPost_uid29_divider_b_1_q_a1_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a10(
	.dataa(!fxp_functions_0_ai8489_a28_sumout),
	.datab(!fxp_functions_0_aMux_121_a1_sumout),
	.datac(!fxp_functions_0_aMux_125_a1_sumout),
	.datad(!fxp_functions_0_aMux_117_a1_sumout),
	.datae(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.dataf(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a10.extended_lut = "off";
defparam fxp_functions_0_ai8489_a10.lut_mask = 64'h555533330F0F00FF;
defparam fxp_functions_0_ai8489_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a11(
	.dataa(!rst),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a4_a_aq),
	.datac(!fxp_functions_0_arShiftCount_uid26_divider_o_a5_a_aq),
	.datad(!fxp_functions_0_aMux_178_a0_combout),
	.datae(!fxp_functions_0_ai8489_a10_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a11.extended_lut = "off";
defparam fxp_functions_0_ai8489_a11.lut_mask = 64'h002080A0002080A0;
defparam fxp_functions_0_ai8489_a11.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai8150_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai8150_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai8150_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai8103_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8103_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8103_a0.extended_lut = "off";
defparam fxp_functions_0_ai8103_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai8103_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a1_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a32_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a1_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_ainvResPostOneHandling2_uid24_divider_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai8126_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0_combout),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq));
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8150_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8150_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8150_a0.extended_lut = "off";
defparam fxp_functions_0_ai8150_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai8150_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8150_a1(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8150_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8150_a1.extended_lut = "off";
defparam fxp_functions_0_ai8150_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai8150_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8150_a2(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8150_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8150_a2.extended_lut = "off";
defparam fxp_functions_0_ai8150_a2.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai8150_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a3_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_wraddr_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_21(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a0_combout),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a1_combout),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a2_combout),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a3_combout),
	.datae(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_cmp_b_a0_a_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_21_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_21.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_21.lut_mask = 64'h0000001000000010;
defparam fxp_functions_0_areduce_nor_21.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai8126_a0(
	.dataa(!rst),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8126_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8126_a0.extended_lut = "off";
defparam fxp_functions_0_ai8126_a0.lut_mask = 64'h8888888888888888;
defparam fxp_functions_0_ai8126_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0.lut_mask = 64'h7575757575757575;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_15_a0(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_15_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_15_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_15_a0.lut_mask = 64'h6666666666666666;
defparam fxp_functions_0_aadd_15_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8126_a1(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8126_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8126_a1.extended_lut = "off";
defparam fxp_functions_0_ai8126_a1.lut_mask = 64'h1EF01EF01EF01EF0;
defparam fxp_functions_0_ai8126_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8126_a2(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8126_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8126_a2.extended_lut = "off";
defparam fxp_functions_0_ai8126_a2.lut_mask = 64'h01FE0FF001FE0FF0;
defparam fxp_functions_0_ai8126_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8126_a3(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq),
	.dataf(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_eq_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8126_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8126_a3.extended_lut = "off";
defparam fxp_functions_0_ai8126_a3.lut_mask = 64'h0001FFFE000FFFF0;
defparam fxp_functions_0_ai8126_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a0(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a1_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a0.extended_lut = "off";
defparam fxp_functions_0_ai6816_a0.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a1(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a6_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a1.extended_lut = "off";
defparam fxp_functions_0_ai6816_a1.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a2(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a11_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a2.extended_lut = "off";
defparam fxp_functions_0_ai6816_a2.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a3(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a16_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a3.extended_lut = "off";
defparam fxp_functions_0_ai6816_a3.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a4(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a21_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a4.extended_lut = "off";
defparam fxp_functions_0_ai6816_a4.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a5(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a26_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a5.extended_lut = "off";
defparam fxp_functions_0_ai6816_a5.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a6(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a31_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a6.extended_lut = "off";
defparam fxp_functions_0_ai6816_a6.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a7(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a36_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a7.extended_lut = "off";
defparam fxp_functions_0_ai6816_a7.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a8(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a41_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a8.extended_lut = "off";
defparam fxp_functions_0_ai6816_a8.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a9(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a46_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a9.extended_lut = "off";
defparam fxp_functions_0_ai6816_a9.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a10(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a51_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a10.extended_lut = "off";
defparam fxp_functions_0_ai6816_a10.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a11(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a56_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a11.extended_lut = "off";
defparam fxp_functions_0_ai6816_a11.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a12(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a61_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a12.extended_lut = "off";
defparam fxp_functions_0_ai6816_a12.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a13(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a66_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a13.extended_lut = "off";
defparam fxp_functions_0_ai6816_a13.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a14(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a71_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a14.extended_lut = "off";
defparam fxp_functions_0_ai6816_a14.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_ai6816_a14.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a15(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a76_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a15.extended_lut = "off";
defparam fxp_functions_0_ai6816_a15.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a15.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a16(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a81_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a16.extended_lut = "off";
defparam fxp_functions_0_ai6816_a16.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a17(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a86_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a17.extended_lut = "off";
defparam fxp_functions_0_ai6816_a17.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a18(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a91_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a18.extended_lut = "off";
defparam fxp_functions_0_ai6816_a18.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a18.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a19(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a96_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a19.extended_lut = "off";
defparam fxp_functions_0_ai6816_a19.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a19.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a20(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a101_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a20.extended_lut = "off";
defparam fxp_functions_0_ai6816_a20.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a20.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a21(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a106_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a21.extended_lut = "off";
defparam fxp_functions_0_ai6816_a21.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a22(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a111_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a22.extended_lut = "off";
defparam fxp_functions_0_ai6816_a22.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a23(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a116_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a23.extended_lut = "off";
defparam fxp_functions_0_ai6816_a23.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a23.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a24(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a121_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a24_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a24.extended_lut = "off";
defparam fxp_functions_0_ai6816_a24.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a24.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a25(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a126_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a25_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a25.extended_lut = "off";
defparam fxp_functions_0_ai6816_a25.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a25.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a26(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a131_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a26_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a26.extended_lut = "off";
defparam fxp_functions_0_ai6816_a26.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a26.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a27(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a136_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a27_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a27.extended_lut = "off";
defparam fxp_functions_0_ai6816_a27.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a27.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a28(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a141_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a28_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a28.extended_lut = "off";
defparam fxp_functions_0_ai6816_a28.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a28.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a29(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a146_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a29_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a29.extended_lut = "off";
defparam fxp_functions_0_ai6816_a29.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a29.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a30(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a151_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a30_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a30.extended_lut = "off";
defparam fxp_functions_0_ai6816_a30.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a30.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a31(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a156_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a31_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a31.extended_lut = "off";
defparam fxp_functions_0_ai6816_a31.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a31.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6816_a32(
	.dataa(!fxp_functions_0_aredist18_normYIsOne_uid16_divider_q_23_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aadd_12_a161_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6816_a32_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6816_a32.extended_lut = "off";
defparam fxp_functions_0_ai6816_a32.lut_mask = 64'h2222222222222222;
defparam fxp_functions_0_ai6816_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_10_a1(
	.dataa(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a_aq),
	.datab(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a_aq),
	.datac(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a_aq),
	.datad(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a_aq),
	.datae(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a_aq),
	.dataf(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_10_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_10_a1.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_10_a1.lut_mask = 64'h8FFF000000000000;
defparam fxp_functions_0_areduce_nor_10_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0(
	.dataa(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a3_a_aq),
	.datab(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a2_a_aq),
	.datac(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a_aq),
	.datad(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0.lut_mask = 64'h50D050D050D050D0;
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1(
	.dataa(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a_aq),
	.datab(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a_aq),
	.datac(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a_aq),
	.datad(!fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1.lut_mask = 64'hB030B030B030B030;
defparam fxp_functions_0_arVStage_uid70_zCount_uid9_divider_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_9(
	.dataa(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a5_a_aq),
	.datab(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a4_a_aq),
	.datac(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a6_a_aq),
	.datad(!fxp_functions_0_avStagei_uid56_zCount_uid9_divider_q_a7_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_9_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_9.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_9.lut_mask = 64'h8000800080008000;
defparam fxp_functions_0_areduce_nor_9.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_17(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_rdcnt_i_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_17_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_17.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_17.lut_mask = 64'h0000001000000010;
defparam fxp_functions_0_areduce_nor_17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a1(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq),
	.datad(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a1.extended_lut = "off";
defparam fxp_functions_0_ai3244_a1.lut_mask = 64'h8000800080008000;
defparam fxp_functions_0_ai3244_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a2(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq),
	.datac(!fxp_functions_0_ai3244_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a2.extended_lut = "off";
defparam fxp_functions_0_ai3244_a2.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_ai3244_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a3(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a3_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq),
	.datad(!fxp_functions_0_ai3244_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a3.extended_lut = "off";
defparam fxp_functions_0_ai3244_a3.lut_mask = 64'h0F4F0F4F0F4F0F4F;
defparam fxp_functions_0_ai3244_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a4(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a2_a_aq),
	.datad(!fxp_functions_0_ai3244_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a4.extended_lut = "off";
defparam fxp_functions_0_ai3244_a4.lut_mask = 64'h555D555D555D555D;
defparam fxp_functions_0_ai3244_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a5(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq),
	.datad(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a5.extended_lut = "off";
defparam fxp_functions_0_ai3244_a5.lut_mask = 64'h8000800080008000;
defparam fxp_functions_0_ai3244_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a6(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a_aq),
	.datac(!fxp_functions_0_ai3244_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a6.extended_lut = "off";
defparam fxp_functions_0_ai3244_a6.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_ai3244_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a7(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a5_a_aq),
	.datad(!fxp_functions_0_ai3244_a6_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a7.extended_lut = "off";
defparam fxp_functions_0_ai3244_a7.lut_mask = 64'h555D555D555D555D;
defparam fxp_functions_0_ai3244_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a8(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a10_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a11_a_aq),
	.datac(!fxp_functions_0_ai3244_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a8.extended_lut = "off";
defparam fxp_functions_0_ai3244_a8.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_ai3244_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a9(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a4_a_aq),
	.datad(!fxp_functions_0_ai3244_a8_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a9.extended_lut = "off";
defparam fxp_functions_0_ai3244_a9.lut_mask = 64'h333B333B333B333B;
defparam fxp_functions_0_ai3244_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a10(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a14_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a12_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a6_a_aq),
	.datad(!fxp_functions_0_ai3244_a8_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a10.extended_lut = "off";
defparam fxp_functions_0_ai3244_a10.lut_mask = 64'h555D555D555D555D;
defparam fxp_functions_0_ai3244_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a11(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a15_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a8_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq),
	.datad(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq),
	.datae(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a7_a_aq),
	.dataf(!fxp_functions_0_ai3244_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a11.extended_lut = "off";
defparam fxp_functions_0_ai3244_a11.lut_mask = 64'h555555555555D555;
defparam fxp_functions_0_ai3244_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3244_a12(
	.dataa(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a13_a_aq),
	.datab(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a9_a_aq),
	.datac(!fxp_functions_0_avStagei_uid50_zCount_uid9_divider_q_a1_a_aq),
	.datad(!fxp_functions_0_ai3244_a6_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3244_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3244_a12.extended_lut = "off";
defparam fxp_functions_0_ai3244_a12.lut_mask = 64'h333B333B333B333B;
defparam fxp_functions_0_ai3244_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_8(
	.dataa(!fxp_functions_0_ai3244_a1_combout),
	.datab(!fxp_functions_0_ai3244_a5_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_8_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_8.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_8.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_areduce_nor_8.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a0(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq),
	.datae(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a0.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_7_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a1(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq),
	.datae(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a1.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a1.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_7_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a2(
	.dataa(!fxp_functions_0_areduce_nor_7_a0_combout),
	.datab(!fxp_functions_0_areduce_nor_7_a1_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a2.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a2.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_areduce_nor_7_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a3(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq),
	.datae(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a3.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a3.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_7_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a4(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq),
	.datae(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a4.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a4.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_7_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7_a5(
	.dataa(!fxp_functions_0_areduce_nor_7_a3_combout),
	.datab(!fxp_functions_0_areduce_nor_7_a4_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7_a5.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7_a5.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_areduce_nor_7_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_7(
	.dataa(!fxp_functions_0_areduce_nor_7_a2_combout),
	.datab(!fxp_functions_0_areduce_nor_7_a5_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_7_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_7.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_7.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_areduce_nor_7.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai1731_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a(
	.clk(clk),
	.d(fxp_functions_0_ai1731_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a(
	.clk(clk),
	.d(fxp_functions_0_ai1731_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai1590_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1590_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1590_a0.extended_lut = "off";
defparam fxp_functions_0_ai1590_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai1590_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a30_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a31_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_inputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq));
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai3159_a1(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a1.extended_lut = "off";
defparam fxp_functions_0_ai3159_a1.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a2(
	.dataa(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a3_a_aq),
	.datab(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq),
	.datae(!fxp_functions_0_ai3159_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a2.extended_lut = "off";
defparam fxp_functions_0_ai3159_a2.lut_mask = 64'h33FF73FF33FF73FF;
defparam fxp_functions_0_ai3159_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a3(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq),
	.datae(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a10_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a3.extended_lut = "off";
defparam fxp_functions_0_ai3159_a3.lut_mask = 64'h0000800000008000;
defparam fxp_functions_0_ai3159_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a4(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq),
	.datac(!fxp_functions_0_areduce_nor_7_a1_combout),
	.datad(!fxp_functions_0_ai3159_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a4.extended_lut = "off";
defparam fxp_functions_0_ai3159_a4.lut_mask = 64'h7777777F7777777F;
defparam fxp_functions_0_ai3159_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a5(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a0_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a5.extended_lut = "off";
defparam fxp_functions_0_ai3159_a5.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a6(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a11_a_aq),
	.datae(!fxp_functions_0_ai3159_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a6.extended_lut = "off";
defparam fxp_functions_0_ai3159_a6.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a7(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a26_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a16_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a1_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a7.extended_lut = "off";
defparam fxp_functions_0_ai3159_a7.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a8(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a14_a_aq),
	.datae(!fxp_functions_0_ai3159_a7_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a8.extended_lut = "off";
defparam fxp_functions_0_ai3159_a8.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a9(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a0_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a9.extended_lut = "off";
defparam fxp_functions_0_ai3159_a9.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a10(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a12_a_aq),
	.datae(!fxp_functions_0_ai3159_a9_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a10.extended_lut = "off";
defparam fxp_functions_0_ai3159_a10.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a11(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a31_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a30_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a15_a_aq),
	.datae(!fxp_functions_0_ai3159_a7_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a11.extended_lut = "off";
defparam fxp_functions_0_ai3159_a11.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a12(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a4_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a12.extended_lut = "off";
defparam fxp_functions_0_ai3159_a12.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a13(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a8_a_aq),
	.datae(!fxp_functions_0_ai3159_a12_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a13.extended_lut = "off";
defparam fxp_functions_0_ai3159_a13.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a14(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a29_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a28_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a13_a_aq),
	.datae(!fxp_functions_0_ai3159_a9_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a14.extended_lut = "off";
defparam fxp_functions_0_ai3159_a14.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a14.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a15(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a27_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a25_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a9_a_aq),
	.datae(!fxp_functions_0_ai3159_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a15.extended_lut = "off";
defparam fxp_functions_0_ai3159_a15.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a15.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a16(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a2_a_aq),
	.datae(!fxp_functions_0_ai3159_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a16.extended_lut = "off";
defparam fxp_functions_0_ai3159_a16.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a17(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a18_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a19_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a17.extended_lut = "off";
defparam fxp_functions_0_ai3159_a17.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a18(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a5_a_aq),
	.datae(!fxp_functions_0_ai3159_a17_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a18.extended_lut = "off";
defparam fxp_functions_0_ai3159_a18.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a18.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a19(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a20_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a21_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a4_a_aq),
	.datae(!fxp_functions_0_ai3159_a17_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a19.extended_lut = "off";
defparam fxp_functions_0_ai3159_a19.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a19.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a20(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq),
	.datad(!fxp_functions_0_areduce_nor_7_a4_combout),
	.datae(!fxp_functions_0_areduce_nor_7_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a20.extended_lut = "off";
defparam fxp_functions_0_ai3159_a20.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_ai3159_a20.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a21(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a6_a_aq),
	.datae(!fxp_functions_0_ai3159_a20_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a21.extended_lut = "off";
defparam fxp_functions_0_ai3159_a21.lut_mask = 64'h777777F7777777F7;
defparam fxp_functions_0_ai3159_a21.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a22(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a24_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a23_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a7_a_aq),
	.datae(!fxp_functions_0_ai3159_a12_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a22.extended_lut = "off";
defparam fxp_functions_0_ai3159_a22.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a22.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3159_a23(
	.dataa(!fxp_functions_0_avCount_uid41_zCount_uid9_divider_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a22_a_aq),
	.datac(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a17_a_aq),
	.datad(!fxp_functions_0_aredist22_in_rsrvd_fix_denominator_1_q_a1_a_aq),
	.datae(!fxp_functions_0_ai3159_a20_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3159_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3159_a23.extended_lut = "off";
defparam fxp_functions_0_ai3159_a23.lut_mask = 64'h5F5F5FDF5F5F5FDF;
defparam fxp_functions_0_ai3159_a23.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a0(
	.dataa(!denominator[30]),
	.datab(!denominator[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a0.lut_mask = 64'h8888888888888888;
defparam fxp_functions_0_areduce_nor_6_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a1(
	.dataa(!denominator[3]),
	.datab(!denominator[0]),
	.datac(!denominator[1]),
	.datad(!denominator[2]),
	.datae(!denominator[4]),
	.dataf(!denominator[5]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a1.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a1.lut_mask = 64'h8000000000000000;
defparam fxp_functions_0_areduce_nor_6_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a2(
	.dataa(!denominator[6]),
	.datab(!denominator[7]),
	.datac(!denominator[8]),
	.datad(!denominator[9]),
	.datae(!denominator[10]),
	.dataf(!denominator[11]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a2.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a2.lut_mask = 64'h8000000000000000;
defparam fxp_functions_0_areduce_nor_6_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a3(
	.dataa(!denominator[12]),
	.datab(!denominator[13]),
	.datac(!denominator[14]),
	.datad(!denominator[15]),
	.datae(!denominator[16]),
	.dataf(!denominator[17]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a3.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a3.lut_mask = 64'h8000000000000000;
defparam fxp_functions_0_areduce_nor_6_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a4(
	.dataa(!denominator[18]),
	.datab(!denominator[19]),
	.datac(!denominator[20]),
	.datad(!denominator[21]),
	.datae(!denominator[22]),
	.dataf(!denominator[23]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a4.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a4.lut_mask = 64'h8000000000000000;
defparam fxp_functions_0_areduce_nor_6_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6_a5(
	.dataa(!denominator[24]),
	.datab(!denominator[25]),
	.datac(!denominator[26]),
	.datad(!denominator[27]),
	.datae(!denominator[28]),
	.dataf(!denominator[29]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6_a5.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6_a5.lut_mask = 64'h8000000000000000;
defparam fxp_functions_0_areduce_nor_6_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_6(
	.dataa(!fxp_functions_0_areduce_nor_6_a0_combout),
	.datab(!fxp_functions_0_areduce_nor_6_a1_combout),
	.datac(!fxp_functions_0_areduce_nor_6_a2_combout),
	.datad(!fxp_functions_0_areduce_nor_6_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_6_a4_combout),
	.dataf(!fxp_functions_0_areduce_nor_6_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_6_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_6.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_6.lut_mask = 64'h0000000000000001;
defparam fxp_functions_0_areduce_nor_6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai1731_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1731_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1731_a0.extended_lut = "off";
defparam fxp_functions_0_ai1731_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai1731_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai1731_a1(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1731_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1731_a1.extended_lut = "off";
defparam fxp_functions_0_ai1731_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai1731_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai1731_a2(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1731_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1731_a2.extended_lut = "off";
defparam fxp_functions_0_ai1731_a2.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai1731_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a3_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_wraddr_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_19(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a2_combout),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a0_combout),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a1_combout),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a3_combout),
	.datae(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_cmp_b_a0_a_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_19_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_19.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_19.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_areduce_nor_19.shared_arith = "off";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a9_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a10_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a11_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a12_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a13_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a0(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a0.lut_mask = 64'h6969696969696969;
defparam fxp_functions_0_aadd_0_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a1(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_0_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a1.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a1.lut_mask = 64'h1E871E871E871E87;
defparam fxp_functions_0_aadd_0_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a2(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_0_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a2.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a2.lut_mask = 64'h01FE7F8001FE7F80;
defparam fxp_functions_0_aadd_0_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_0_a3(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq),
	.dataf(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_eq_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_0_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_0_a3.extended_lut = "off";
defparam fxp_functions_0_aadd_0_a3.lut_mask = 64'h0001FFFE007FFF80;
defparam fxp_functions_0_aadd_0_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a8_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_2(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a3_a_aq),
	.datae(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_2_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_2.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_2.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_areduce_nor_2.shared_arith = "off";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist8_lowRangeB_uid98_invPolyEval_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a23_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a24_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a25_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a26_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a27_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a28_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_as2sumAHighB_uid100_invPolyEval_o_a29_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai6157_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai6102_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6102_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6102_a0.extended_lut = "off";
defparam fxp_functions_0_ai6102_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai6102_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_inputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a7_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6157_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6157_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6157_a0.extended_lut = "off";
defparam fxp_functions_0_ai6157_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai6157_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_13(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a0_combout),
	.datae(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_13_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_13.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_13.lut_mask = 64'h000000D8000000D8;
defparam fxp_functions_0_areduce_nor_13.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a6_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai6114_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6114_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6114_a0.extended_lut = "off";
defparam fxp_functions_0_ai6114_a0.lut_mask = 64'h6363636363636363;
defparam fxp_functions_0_ai6114_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6114_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6114_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6114_a1.extended_lut = "off";
defparam fxp_functions_0_ai6114_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fxp_functions_0_ai6114_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai6114_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq),
	.datae(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai6114_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai6114_a2.extended_lut = "off";
defparam fxp_functions_0_ai6114_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fxp_functions_0_ai6114_a2.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a5_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a28_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a28_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a29_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a29_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a30_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a30_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a31_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a31_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a32_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a32_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a33_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a33_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a34_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a34_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a35_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a35_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a36_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a36_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a37_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a37_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a38_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a38_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a39_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a39_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a40_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a40_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a41_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a41_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a42_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a42_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_s0_a43_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_delay_adelay_signals_a0_a_a43_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_14(
	.dataa(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist2_yAddr_uid19_divider_merged_bit_select_b_22_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_14_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_14.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_14.lut_mask = 64'h1010101010101010;
defparam fxp_functions_0_areduce_nor_14.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a4_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a(
	.clk(clk),
	.d(fxp_functions_0_ai3830_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a(
	.clk(clk),
	.d(fxp_functions_0_ai3830_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai1992_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1992_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1992_a0.extended_lut = "off";
defparam fxp_functions_0_ai1992_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai1992_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist9_lowRangeB_uid92_invPolyEval_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_as1sumAHighB_uid94_invPolyEval_o_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ch_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_outputreg0_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid112_pT2_uid97_invPolyEval_cma_ah_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_inputreg0_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a3_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai3830_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3830_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3830_a0.extended_lut = "off";
defparam fxp_functions_0_ai3830_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai3830_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3830_a1(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3830_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3830_a1.extended_lut = "off";
defparam fxp_functions_0_ai3830_a1.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai3830_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_cmp_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_20(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_wraddr_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq),
	.datae(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_20_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_20.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_20.lut_mask = 64'h08085D0808085D08;
defparam fxp_functions_0_areduce_nor_20.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a2_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im10_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai1997_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai1997_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai1997_a0.extended_lut = "off";
defparam fxp_functions_0_ai1997_a0.lut_mask = 64'h6666666666666666;
defparam fxp_functions_0_ai1997_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aadd_2_a0(
	.dataa(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist5_yAddr_uid19_divider_merged_bit_select_c_17_rdcnt_i_a1_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aadd_2_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aadd_2_a0.extended_lut = "off";
defparam fxp_functions_0_aadd_2_a0.lut_mask = 64'h6666666666666666;
defparam fxp_functions_0_aadd_2_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a14_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a1_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a15_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a16_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a17_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a19_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a20_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a21_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a22_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a22_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a23_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a23_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a24_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a24_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a25_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a25_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a26_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a26_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a(
	.clk(clk),
	.d(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_s0_a27_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_delay_adelay_signals_a0_a_a27_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_ff fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_s0_a0_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a_aq));
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a(
	.clk(clk),
	.d(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_s0_a18_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a_aq));
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_delay_adelay_signals_a0_a_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist6_memoryC3_uid83_invTabGen_lutmem_r_1_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ch_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.sclr1(gnd),
	.q(fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a_aq));
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aprodXY_uid109_pT1_uid91_invPolyEval_cma_ah_a0_a_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai3634_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai2020_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai2020_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai2020_a0.extended_lut = "off";
defparam fxp_functions_0_ai2020_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai2020_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a8_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a8_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a9_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a9_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a10_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a10_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a11_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a11_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a12_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a12_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a13_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a13_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a14_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a14_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a15_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a15_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a16_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a16_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a17_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a17_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a18_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a18_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a19_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a19_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a20_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a20_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a21_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a21_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a22_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a22_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai3634_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai3634_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai3634_a0.extended_lut = "off";
defparam fxp_functions_0_ai3634_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai3634_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_4(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a0_combout),
	.datae(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_4_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_4.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_4.lut_mask = 64'h000000D8000000D8;
defparam fxp_functions_0_areduce_nor_4.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist3_yAddr_uid19_divider_merged_bit_select_c_3_q_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a.extended_lut = "off";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_enaAnd_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai2032_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai2032_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai2032_a0.extended_lut = "off";
defparam fxp_functions_0_ai2032_a0.lut_mask = 64'h6363636363636363;
defparam fxp_functions_0_ai2032_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai2032_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai2032_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai2032_a1.extended_lut = "off";
defparam fxp_functions_0_ai2032_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fxp_functions_0_ai2032_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai2032_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datae(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai2032_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai2032_a2.extended_lut = "off";
defparam fxp_functions_0_ai2032_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fxp_functions_0_ai2032_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_8_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_8_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_8_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_8_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_8_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_16_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_16_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_16_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_16_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_16_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_12_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_12_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_12_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_12_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_12_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_20_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_20_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_20_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_20_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_20_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_10_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_10_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_10_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_10_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_10_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_18_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_18_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_18_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_18_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_18_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_14_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_14_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_14_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_14_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_14_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_22_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_22_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_22_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_22_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_22_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_9_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_9_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_9_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_9_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_9_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_17_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_17_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_17_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_17_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_17_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_13_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_13_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_13_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_13_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_13_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_21_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_21_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_21_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_21_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_21_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_11_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_11_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_11_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_11_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_11_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_19_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_19_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_19_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_19_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_19_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_15_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_15_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_15_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_15_a1.lut_mask = 64'h048C048C048C048C;
defparam fxp_functions_0_aMux_15_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_23_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_23_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_23_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_23_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_23_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a0.lut_mask = 64'h0020002000200020;
defparam fxp_functions_0_aMux_40_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a1.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_40_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_19_a0_combout),
	.datad(!fxp_functions_0_aMux_11_a1_combout),
	.datae(!fxp_functions_0_aMux_40_a0_combout),
	.dataf(!fxp_functions_0_aMux_40_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a2.lut_mask = 64'h0123CDEFCDEFCDEF;
defparam fxp_functions_0_aMux_40_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a3(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a3.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a3.lut_mask = 64'h0020002000200020;
defparam fxp_functions_0_aMux_40_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a4(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a4.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a4.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_40_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a5(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_18_a0_combout),
	.datad(!fxp_functions_0_aMux_10_a1_combout),
	.datae(!fxp_functions_0_aMux_40_a3_combout),
	.dataf(!fxp_functions_0_aMux_40_a4_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a5.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a5.lut_mask = 64'h0123CDEFCDEFCDEF;
defparam fxp_functions_0_aMux_40_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a6(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a6.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a6.lut_mask = 64'h0020002000200020;
defparam fxp_functions_0_aMux_40_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a7(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a7.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a7.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_40_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a8(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_17_a0_combout),
	.datad(!fxp_functions_0_aMux_9_a1_combout),
	.datae(!fxp_functions_0_aMux_40_a6_combout),
	.dataf(!fxp_functions_0_aMux_40_a7_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a8.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a8.lut_mask = 64'h0123CDEFCDEFCDEF;
defparam fxp_functions_0_aMux_40_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_32_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_32_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_32_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_32_a0.lut_mask = 64'h0020002000200020;
defparam fxp_functions_0_aMux_32_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_32_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_32_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_32_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_32_a1.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_32_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a9(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_16_a0_combout),
	.datad(!fxp_functions_0_aMux_8_a1_combout),
	.datae(!fxp_functions_0_aMux_32_a0_combout),
	.dataf(!fxp_functions_0_aMux_32_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a9.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a9.lut_mask = 64'h0123CDEFCDEFCDEF;
defparam fxp_functions_0_aMux_40_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a10(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a10.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a10.lut_mask = 64'h2020202020202020;
defparam fxp_functions_0_aMux_40_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a11(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a11.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a11.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_40_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a12(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq),
	.datad(!fxp_functions_0_aMux_40_a10_combout),
	.datae(!fxp_functions_0_aMux_40_a1_combout),
	.dataf(!fxp_functions_0_aMux_40_a11_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a12.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a12.lut_mask = 64'h00275577AAAFFFFF;
defparam fxp_functions_0_aMux_40_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a13(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a_aq),
	.dataf(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a13.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a13.lut_mask = 64'h001040508090C0D0;
defparam fxp_functions_0_aMux_40_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a14(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq),
	.datad(!fxp_functions_0_aMux_40_a10_combout),
	.datae(!fxp_functions_0_aMux_40_a4_combout),
	.dataf(!fxp_functions_0_aMux_40_a13_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a14.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a14.lut_mask = 64'h00275577AAAFFFFF;
defparam fxp_functions_0_aMux_40_a14.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a15(
	.dataa(!fxp_functions_0_aMux_40_a6_combout),
	.datab(!fxp_functions_0_aMux_40_a7_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a15.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a15.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aMux_40_a15.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a16(
	.dataa(!fxp_functions_0_aMux_40_a0_combout),
	.datab(!fxp_functions_0_aMux_40_a1_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a16.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a16.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aMux_40_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_72_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aMux_64_a6_combout),
	.datad(!fxp_functions_0_aMux_40_a9_combout),
	.datae(!fxp_functions_0_aMux_40_a14_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_72_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_72_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_72_a0.lut_mask = 64'h0C1D2E3F0C1D2E3F;
defparam fxp_functions_0_aMux_72_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a(
	.clk(clk),
	.d(fxp_functions_0_ai4289_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a2_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a0_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_ardaddr_reg_a2_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_ai4258_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_sticky_ena_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_cmpReg_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai4258_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai4258_a0.extended_lut = "off";
defparam fxp_functions_0_ai4258_a0.lut_mask = 64'h3737373737373737;
defparam fxp_functions_0_ai4258_a0.shared_arith = "off";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a7_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a1_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a12_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a2_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a17_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a3_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a22_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a4_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a27_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a5_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a32_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a6_a.power_up = "dont_care";

fourteennm_ff fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a(
	.clk(clk),
	.d(fxp_functions_0_aMux_72_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a_aq));
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.is_wysiwyg = "true";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_mem_dmem_aauto_generated_aaltera_syncram_impl1_aportadatain_reg_a7_a.power_up = "dont_care";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_5(
	.dataa(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist4_yAddr_uid19_divider_merged_bit_select_c_10_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_5_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_5.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_5.lut_mask = 64'h1010101010101010;
defparam fxp_functions_0_areduce_nor_5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_30_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_30_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_30_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_30_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_30_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_26_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_26_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_26_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_26_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_26_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_54_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_22_a0_combout),
	.datad(!fxp_functions_0_aMux_30_a0_combout),
	.datae(!fxp_functions_0_aMux_26_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_54_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_54_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_54_a0.lut_mask = 64'h084C2A6E084C2A6E;
defparam fxp_functions_0_aMux_54_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_94_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_94_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_94_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_94_a1.lut_mask = 64'h8080808080808080;
defparam fxp_functions_0_aMux_94_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_56_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.datad(!fxp_functions_0_aMux_94_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_56_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_56_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_56_a1.lut_mask = 64'h0027002700270027;
defparam fxp_functions_0_aMux_56_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_31_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_31_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_31_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_31_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_31_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_27_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_27_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_27_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_27_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_27_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_55_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_23_a0_combout),
	.datad(!fxp_functions_0_aMux_31_a0_combout),
	.datae(!fxp_functions_0_aMux_27_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_55_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_55_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_55_a0.lut_mask = 64'h084C2A6E084C2A6E;
defparam fxp_functions_0_aMux_55_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_57_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.datad(!fxp_functions_0_aMux_94_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_57_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_57_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_57_a1.lut_mask = 64'h0027002700270027;
defparam fxp_functions_0_aMux_57_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_29_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_29_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_29_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_29_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_29_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_25_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_25_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_25_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_25_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_25_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_53_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_21_a0_combout),
	.datad(!fxp_functions_0_aMux_29_a0_combout),
	.datae(!fxp_functions_0_aMux_25_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_53_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_53_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_53_a0.lut_mask = 64'h084C2A6E084C2A6E;
defparam fxp_functions_0_aMux_53_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_28_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_28_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_28_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_28_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_28_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_24_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_24_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_24_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_24_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_24_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_52_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aMux_20_a0_combout),
	.datad(!fxp_functions_0_aMux_28_a0_combout),
	.datae(!fxp_functions_0_aMux_24_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_52_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_52_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_52_a0.lut_mask = 64'h084C2A6E084C2A6E;
defparam fxp_functions_0_aMux_52_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai4289_a0(
	.dataa(!rst),
	.datab(!en[0]),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai4289_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai4289_a0.extended_lut = "off";
defparam fxp_functions_0_ai4289_a0.lut_mask = 64'h5D7F5D7F5D7F5D7F;
defparam fxp_functions_0_ai4289_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2.lut_mask = 64'h2727272727272727;
defparam fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_11(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_wraddr_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datad(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a0_combout),
	.datae(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdmux_q_a0_a_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_11_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_11.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_11.lut_mask = 64'h000000D8000000D8;
defparam fxp_functions_0_areduce_nor_11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_63_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_63_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_63_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_63_a0.lut_mask = 64'h0000800000008000;
defparam fxp_functions_0_aMux_63_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_61_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_61_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_61_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_61_a0.lut_mask = 64'h0000800000008000;
defparam fxp_functions_0_aMux_61_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_62_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_62_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_62_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_62_a0.lut_mask = 64'h0000800000008000;
defparam fxp_functions_0_aMux_62_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_93_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aMux_63_a0_combout),
	.datad(!fxp_functions_0_aMux_61_a0_combout),
	.datae(!fxp_functions_0_aMux_62_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_93_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_93_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_93_a0.lut_mask = 64'h048C26AE048C26AE;
defparam fxp_functions_0_aMux_93_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_60_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a4_a_aq),
	.datad(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a5_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_60_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_60_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_60_a0.lut_mask = 64'h0000800000008000;
defparam fxp_functions_0_aMux_60_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_59_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.datad(!fxp_functions_0_aMux_94_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_59_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_59_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_59_a1.lut_mask = 64'h0027002700270027;
defparam fxp_functions_0_aMux_59_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_58_a1(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datad(!fxp_functions_0_aMux_94_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_58_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_58_a1.extended_lut = "off";
defparam fxp_functions_0_aMux_58_a1.lut_mask = 64'h0027002700270027;
defparam fxp_functions_0_aMux_58_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai4270_a0(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai4270_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai4270_a0.extended_lut = "off";
defparam fxp_functions_0_ai4270_a0.lut_mask = 64'h6363636363636363;
defparam fxp_functions_0_ai4270_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai4270_a1(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai4270_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai4270_a1.extended_lut = "off";
defparam fxp_functions_0_ai4270_a1.lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam fxp_functions_0_ai4270_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai4270_a2(
	.dataa(!en[0]),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datad(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datae(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_eq_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai4270_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai4270_a2.extended_lut = "off";
defparam fxp_functions_0_ai4270_a2.lut_mask = 64'h01FE55AA01FE55AA;
defparam fxp_functions_0_ai4270_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_95_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aMux_63_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_95_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_95_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_95_a0.lut_mask = 64'h0808080808080808;
defparam fxp_functions_0_aMux_95_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_94_a2(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datac(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a2_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.dataf(!fxp_functions_0_aMux_94_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_94_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_94_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_94_a2.lut_mask = 64'h00000000008020A0;
defparam fxp_functions_0_aMux_94_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_12(
	.dataa(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a0_a_aq),
	.datab(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a1_a_aq),
	.datac(!fxp_functions_0_aredist0_yAddr_uid19_divider_merged_bit_select_b_7_rdcnt_i_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_12_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_12.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_12.lut_mask = 64'h1010101010101010;
defparam fxp_functions_0_areduce_nor_12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a17_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a18_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a19_a_aq),
	.datad(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a20_a_aq),
	.datae(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a21_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a22_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a6_a_aq),
	.datad(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a7_a_aq),
	.datae(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a8_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a10_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a11_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a12_a_aq),
	.datad(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a13_a_aq),
	.datae(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a14_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a16_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a3_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a24_a_aq),
	.datad(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a23_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4.lut_mask = 64'h8000800080008000;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a28_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a30_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a29_a_aq),
	.datad(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a27_a_aq),
	.datae(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a26_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a4_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a5_a_aq),
	.datac(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a25_a_aq),
	.datad(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a4_combout),
	.datae(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a9_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a15_a_aq),
	.datac(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a2_combout),
	.datad(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a3_combout),
	.datae(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a6_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7.lut_mask = 64'h0000000800000008;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0(
	.dataa(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist20_normYNoLeadOne_uid11_divider_b_1_q_a1_a_aq),
	.datac(!fxp_functions_0_aredist19_normYIsOneC2_uid15_divider_b_1_q_a0_a_aq),
	.datad(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a1_combout),
	.datae(!fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a7_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0.lut_mask = 64'h0000000800000008;
defparam fxp_functions_0_anormYIsOne_uid16_divider_qi_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_32_a2(
	.dataa(!fxp_functions_0_aMux_32_a0_combout),
	.datab(!fxp_functions_0_aMux_32_a1_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_32_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_32_a2.extended_lut = "off";
defparam fxp_functions_0_aMux_32_a2.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aMux_32_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_40_a17(
	.dataa(!fxp_functions_0_aMux_40_a3_combout),
	.datab(!fxp_functions_0_aMux_40_a4_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_40_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_40_a17.extended_lut = "off";
defparam fxp_functions_0_aMux_40_a17.lut_mask = 64'h7777777777777777;
defparam fxp_functions_0_aMux_40_a17.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aMux_64_a0(
	.dataa(!fxp_functions_0_aredist10_r_uid72_zCount_uid9_divider_q_1_q_a0_a_aq),
	.datab(!fxp_functions_0_aMux_64_a6_combout),
	.datac(!fxp_functions_0_aMux_64_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aMux_64_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aMux_64_a0.extended_lut = "off";
defparam fxp_functions_0_aMux_64_a0.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fxp_functions_0_aMux_64_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a0(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a7_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a23_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a15_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a27_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a28_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a0.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a0.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_18_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a1(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a19_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a18_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a10_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a4_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a20_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a1.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a1.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_18_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a2(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a0_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a16_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a8_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a24_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a25_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a2.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a2.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_18_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a3(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a1_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a17_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a9_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a22_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a3.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a3.lut_mask = 64'h8000800080008000;
defparam fxp_functions_0_areduce_nor_18_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a4(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a3_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a11_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a5_a_aq),
	.datad(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a21_a_aq),
	.datae(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a4.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a4.lut_mask = 64'h8000000080000000;
defparam fxp_functions_0_areduce_nor_18_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a5(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a13_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a6_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a14_a_aq),
	.datad(!fxp_functions_0_areduce_nor_18_a3_combout),
	.datae(!fxp_functions_0_areduce_nor_18_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a5.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a5.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_areduce_nor_18_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18_a6(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a12_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a26_a_aq),
	.datac(!fxp_functions_0_areduce_nor_18_a1_combout),
	.datad(!fxp_functions_0_areduce_nor_18_a2_combout),
	.datae(!fxp_functions_0_areduce_nor_18_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18_a6.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18_a6.lut_mask = 64'h0000000800000008;
defparam fxp_functions_0_areduce_nor_18_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_areduce_nor_18(
	.dataa(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a29_a_aq),
	.datab(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a30_a_aq),
	.datac(!fxp_functions_0_aredist23_in_rsrvd_fix_denominator_4_q_a31_a_aq),
	.datad(!fxp_functions_0_areduce_nor_18_a0_combout),
	.datae(!fxp_functions_0_areduce_nor_18_a6_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_areduce_nor_18_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_areduce_nor_18.extended_lut = "off";
defparam fxp_functions_0_areduce_nor_18.lut_mask = 64'h0000008000000080;
defparam fxp_functions_0_areduce_nor_18.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a32(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_109_a1_sumout),
	.datad(!fxp_functions_0_aMux_105_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a32_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a32.extended_lut = "off";
defparam fxp_functions_0_ai8489_a32.lut_mask = 64'h8C9D8C9D8C9D8C9D;
defparam fxp_functions_0_ai8489_a32.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_ai8489_a33(
	.dataa(!fxp_functions_0_arShiftCount_uid26_divider_o_a3_a_aq),
	.datab(!fxp_functions_0_arShiftCount_uid26_divider_o_a2_a_aq),
	.datac(!fxp_functions_0_aMux_104_a1_sumout),
	.datad(!fxp_functions_0_aMux_108_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_ai8489_a33_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_ai8489_a33.extended_lut = "off";
defparam fxp_functions_0_ai8489_a33.lut_mask = 64'h89CD89CD89CD89CD;
defparam fxp_functions_0_ai8489_a33.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0.extended_lut = "off";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ch_a0_a_a14_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0.extended_lut = "off";
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_aprodXInvY_uid27_divider_im0_cma_ah_a0_a_a15_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0.extended_lut = "off";
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_aprodXInvY_uid27_divider_ma5_cma_ah_a0_a_a14_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ch_a1_a_a17_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a1_a_a1.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a2_a_a2.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a3_a_a3.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a1_a_a4_a_a4.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a1_a_a6.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a2_a_a7.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a3_a_a8.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a4_a_a9.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a5_a_a10.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a6_a_a11.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a7_a_a12.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a8_a_a13.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a9_a_a14.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a10_a_a15.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16.extended_lut = "off";
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_amultSumOfTwoTS_uid142_pT3_uid103_invPolyEval_cma_ah_a0_a_a11_a_a16.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0.extended_lut = "off";
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0.lut_mask = 64'h0000000000000000;
defparam fxp_functions_0_asm0_uid141_pT3_uid103_invPolyEval_cma_ah_a0_a_a17_a_a0.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a0_a_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a1_a_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a2_a_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a3_a_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist11_r_uid72_zCount_uid9_divider_q_32_outputreg0_q_a4_a_a_wirecell.shared_arith = "off";

fourteennm_lcell_comb fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell(
	.dataa(!fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_aq),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell.extended_lut = "off";
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fxp_functions_0_aredist21_in_rsrvd_fix_numerator_29_rdcnt_i_a0_a_a_wirecell.shared_arith = "off";

assign result[0] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a0_combout;

assign result[10] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a10_combout;

assign result[11] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a11_combout;

assign result[12] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a12_combout;

assign result[13] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a13_combout;

assign result[14] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a14_combout;

assign result[15] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a15_combout;

assign result[16] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a16_combout;

assign result[17] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a17_combout;

assign result[18] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a18_combout;

assign result[19] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a19_combout;

assign result[1] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a1_combout;

assign result[20] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a20_combout;

assign result[21] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a21_combout;

assign result[22] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a22_combout;

assign result[23] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a23_combout;

assign result[24] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a24_combout;

assign result[25] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a25_combout;

assign result[26] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a26_combout;

assign result[27] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a27_combout;

assign result[28] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a28_combout;

assign result[29] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a29_combout;

assign result[2] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a2_combout;

assign result[30] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a30_combout;

assign result[31] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a31_combout;

assign result[3] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a3_combout;

assign result[4] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a4_combout;

assign result[5] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a5_combout;

assign result[6] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a6_combout;

assign result[7] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a7_combout;

assign result[8] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a8_combout;

assign result[9] = fxp_functions_0_aresFinal_uid37_divider_q_a0_a_a9_combout;

endmodule
