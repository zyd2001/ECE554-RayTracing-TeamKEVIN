module mem_main_scalar_test();


endmodule