module IC();



endmodule