module IC();

endmodule