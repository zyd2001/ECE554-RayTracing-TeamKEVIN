// Fix_Sqrt.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module Fix_Sqrt (
		input  wire        clk,     //     clk.clk
		input  wire        rst,     //     rst.reset
		input  wire [0:0]  en,      //      en.en
		input  wire [31:0] radical, // radical.radical
		output wire [31:0] result   //  result.result
	);

	Fix_Sqrt_altera_fxp_functions_191_pjm2y2i fxp_functions_0 (
		.clk     (clk),     //   input,   width = 1,     clk.clk
		.rst     (rst),     //   input,   width = 1,     rst.reset
		.en      (en),      //   input,   width = 1,      en.en
		.radical (radical), //   input,  width = 32, radical.radical
		.result  (result)   //  output,  width = 32,  result.result
	);

endmodule
