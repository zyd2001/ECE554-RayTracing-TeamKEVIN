// FPU.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module FPU (
		input  wire        clk,       // s1.clk
		input  wire        clk_en,    //   .clk_en
		input  wire [31:0] dataa,     //   .dataa
		input  wire [31:0] datab,     //   .datab
		input  wire [2:0]  n,         //   .n
		input  wire        reset,     //   .reset
		input  wire        reset_req, //   .reset_req
		input  wire        start,     //   .start
		output wire        done,      //   .done
		output wire [31:0] result     //   .result
	);

	fpoint2_multi #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1)
	) nios_custom_instr_floating_point_2_multi_0 (
		.clk       (clk),       //   input,   width = 1, s1.clk
		.clk_en    (clk_en),    //   input,   width = 1,   .clk_en
		.dataa     (dataa),     //   input,  width = 32,   .dataa
		.datab     (datab),     //   input,  width = 32,   .datab
		.n         (n),         //   input,   width = 3,   .n
		.reset     (reset),     //   input,   width = 1,   .reset
		.reset_req (reset_req), //   input,   width = 1,   .reset_req
		.start     (start),     //   input,   width = 1,   .start
		.done      (done),      //  output,   width = 1,   .done
		.result    (result)     //  output,  width = 32,   .result
	);

endmodule
